package global_package;


// Constants

localparam bit unsigned [639:0] FINAL_PAD = 640'h8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000580;

localparam bit unsigned [1023:0] IPAD = 1024'h3636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636363636;

localparam bit unsigned [1023:0] OPAD = 1024'h5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C;


// Functions

function bit unsigned [1023:0] hmac_padded(bit unsigned [383:0] hmac_digest);
  return ((hmac_digest << 384'd640) | FINAL_PAD);
endfunction

function bit unsigned [1023:0] key_ipadded(bit unsigned [383:0] key);
  return ((key << 384'd640) ^ IPAD);
endfunction

function bit unsigned [1023:0] key_opadded(bit unsigned [383:0] key);
  return ((key << 384'd640) ^ OPAD);
endfunction


endpackage
