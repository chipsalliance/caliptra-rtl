//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
// DESCRIPTION: Base sequence to perform a mailbox command within the
//              soc_ifc environment.
//              Extended to provide additional functionality.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
class soc_ifc_env_axi_uvm_b2b_rand_sequence extends aaxi_uvm_seq_base; //soc_ifc_env_sequence_base #(.CONFIG_T(soc_ifc_env_configuration_t));


    `uvm_object_utils( soc_ifc_env_axi_uvm_b2b_rand_sequence )
  
    uvm_status_e reg_sts;

    extern virtual task read_reg();
    extern virtual task write_reg(int id);
    extern virtual task read_write_reg(int id);

    function new(string name = "");
        super.new(name);
    endfunction

    virtual task pre_body();
        super.pre_body();
    endtask

    virtual task body();
        write_reg(0);
        read_reg();
        #1000ns;
        read_write_reg('h0);
    endtask
  
endclass

task soc_ifc_env_axi_uvm_b2b_rand_sequence::read_reg();
endtask

task soc_ifc_env_axi_uvm_b2b_rand_sequence::write_reg(int id);
endtask

task soc_ifc_env_axi_uvm_b2b_rand_sequence::read_write_reg(int id);
endtask
