// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef CALIPTRA_REG_DEFINES_HEADER
`define CALIPTRA_REG_DEFINES_HEADER


`define CLP_BASE_ADDR                                                                               (32'h0)
`define CLP_DOE_REG_BASE_ADDR                                                                       (32'h10000000)
`define CLP_DOE_REG_DOE_IV_0                                                                        (32'h10000000)
`define DOE_REG_DOE_IV_0                                                                            (32'h0)
`define CLP_DOE_REG_DOE_IV_1                                                                        (32'h10000004)
`define DOE_REG_DOE_IV_1                                                                            (32'h4)
`define CLP_DOE_REG_DOE_IV_2                                                                        (32'h10000008)
`define DOE_REG_DOE_IV_2                                                                            (32'h8)
`define CLP_DOE_REG_DOE_IV_3                                                                        (32'h1000000c)
`define DOE_REG_DOE_IV_3                                                                            (32'hc)
`define CLP_DOE_REG_DOE_CTRL                                                                        (32'h10000010)
`define DOE_REG_DOE_CTRL                                                                            (32'h10)
`define DOE_REG_DOE_CTRL_CMD_LOW                                                                    (0)
`define DOE_REG_DOE_CTRL_CMD_MASK                                                                   (32'h3)
`define DOE_REG_DOE_CTRL_DEST_LOW                                                                   (2)
`define DOE_REG_DOE_CTRL_DEST_MASK                                                                  (32'h7c)
`define CLP_DOE_REG_DOE_STATUS                                                                      (32'h10000014)
`define DOE_REG_DOE_STATUS                                                                          (32'h14)
`define DOE_REG_DOE_STATUS_READY_LOW                                                                (0)
`define DOE_REG_DOE_STATUS_READY_MASK                                                               (32'h1)
`define DOE_REG_DOE_STATUS_VALID_LOW                                                                (1)
`define DOE_REG_DOE_STATUS_VALID_MASK                                                               (32'h2)
`define DOE_REG_DOE_STATUS_UDS_FLOW_DONE_LOW                                                        (2)
`define DOE_REG_DOE_STATUS_UDS_FLOW_DONE_MASK                                                       (32'h4)
`define DOE_REG_DOE_STATUS_FE_FLOW_DONE_LOW                                                         (3)
`define DOE_REG_DOE_STATUS_FE_FLOW_DONE_MASK                                                        (32'h8)
`define DOE_REG_DOE_STATUS_DEOBF_SECRETS_CLEARED_LOW                                                (4)
`define DOE_REG_DOE_STATUS_DEOBF_SECRETS_CLEARED_MASK                                               (32'h10)
`define CLP_DOE_REG_INTR_BLOCK_RF_START                                                             (32'h10000800)
`define CLP_DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10000800)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                      (32'h800)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                         (0)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                        (32'h1)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                         (1)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                        (32'h2)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10000804)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                       (32'h804)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                         (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                        (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                         (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                        (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                         (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                        (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                         (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                        (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10000808)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                       (32'h808)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                 (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                                (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1000080c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                   (32'h80c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10000810)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                   (32'h810)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10000814)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                 (32'h814)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                                  (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                                 (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                                  (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                                 (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                                  (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                                 (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                                  (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                                 (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10000818)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                 (32'h818)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                          (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                         (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1000081c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                     (32'h81c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                     (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                    (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                     (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                    (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                     (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                    (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                     (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                    (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10000820)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                     (32'h820)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                             (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                            (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                               (32'h10000900)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                   (32'h900)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                               (32'h10000904)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                   (32'h904)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                               (32'h10000908)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                   (32'h908)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                               (32'h1000090c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                   (32'h90c)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10000980)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                           (32'h980)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                          (32'h10000a00)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                              (32'ha00)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                          (32'h10000a04)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                              (32'ha04)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                          (32'h10000a08)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                              (32'ha08)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                          (32'h10000a0c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                              (32'ha0c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10000a10)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                      (32'ha10)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_ECC_REG_BASE_ADDR                                                                       (32'h10008000)
`define CLP_ECC_REG_ECC_NAME_0                                                                      (32'h10008000)
`define ECC_REG_ECC_NAME_0                                                                          (32'h0)
`define CLP_ECC_REG_ECC_NAME_1                                                                      (32'h10008004)
`define ECC_REG_ECC_NAME_1                                                                          (32'h4)
`define CLP_ECC_REG_ECC_VERSION_0                                                                   (32'h10008008)
`define ECC_REG_ECC_VERSION_0                                                                       (32'h8)
`define CLP_ECC_REG_ECC_VERSION_1                                                                   (32'h1000800c)
`define ECC_REG_ECC_VERSION_1                                                                       (32'hc)
`define CLP_ECC_REG_ECC_CTRL                                                                        (32'h10008010)
`define ECC_REG_ECC_CTRL                                                                            (32'h10)
`define ECC_REG_ECC_CTRL_CTRL_LOW                                                                   (0)
`define ECC_REG_ECC_CTRL_CTRL_MASK                                                                  (32'h3)
`define ECC_REG_ECC_CTRL_ZEROIZE_LOW                                                                (2)
`define ECC_REG_ECC_CTRL_ZEROIZE_MASK                                                               (32'h4)
`define ECC_REG_ECC_CTRL_PCR_SIGN_LOW                                                               (3)
`define ECC_REG_ECC_CTRL_PCR_SIGN_MASK                                                              (32'h8)
`define ECC_REG_ECC_CTRL_DH_SHAREDKEY_LOW                                                           (4)
`define ECC_REG_ECC_CTRL_DH_SHAREDKEY_MASK                                                          (32'h10)
`define CLP_ECC_REG_ECC_STATUS                                                                      (32'h10008018)
`define ECC_REG_ECC_STATUS                                                                          (32'h18)
`define ECC_REG_ECC_STATUS_READY_LOW                                                                (0)
`define ECC_REG_ECC_STATUS_READY_MASK                                                               (32'h1)
`define ECC_REG_ECC_STATUS_VALID_LOW                                                                (1)
`define ECC_REG_ECC_STATUS_VALID_MASK                                                               (32'h2)
`define CLP_ECC_REG_ECC_SEED_0                                                                      (32'h10008080)
`define ECC_REG_ECC_SEED_0                                                                          (32'h80)
`define CLP_ECC_REG_ECC_SEED_1                                                                      (32'h10008084)
`define ECC_REG_ECC_SEED_1                                                                          (32'h84)
`define CLP_ECC_REG_ECC_SEED_2                                                                      (32'h10008088)
`define ECC_REG_ECC_SEED_2                                                                          (32'h88)
`define CLP_ECC_REG_ECC_SEED_3                                                                      (32'h1000808c)
`define ECC_REG_ECC_SEED_3                                                                          (32'h8c)
`define CLP_ECC_REG_ECC_SEED_4                                                                      (32'h10008090)
`define ECC_REG_ECC_SEED_4                                                                          (32'h90)
`define CLP_ECC_REG_ECC_SEED_5                                                                      (32'h10008094)
`define ECC_REG_ECC_SEED_5                                                                          (32'h94)
`define CLP_ECC_REG_ECC_SEED_6                                                                      (32'h10008098)
`define ECC_REG_ECC_SEED_6                                                                          (32'h98)
`define CLP_ECC_REG_ECC_SEED_7                                                                      (32'h1000809c)
`define ECC_REG_ECC_SEED_7                                                                          (32'h9c)
`define CLP_ECC_REG_ECC_SEED_8                                                                      (32'h100080a0)
`define ECC_REG_ECC_SEED_8                                                                          (32'ha0)
`define CLP_ECC_REG_ECC_SEED_9                                                                      (32'h100080a4)
`define ECC_REG_ECC_SEED_9                                                                          (32'ha4)
`define CLP_ECC_REG_ECC_SEED_10                                                                     (32'h100080a8)
`define ECC_REG_ECC_SEED_10                                                                         (32'ha8)
`define CLP_ECC_REG_ECC_SEED_11                                                                     (32'h100080ac)
`define ECC_REG_ECC_SEED_11                                                                         (32'hac)
`define CLP_ECC_REG_ECC_MSG_0                                                                       (32'h10008100)
`define ECC_REG_ECC_MSG_0                                                                           (32'h100)
`define CLP_ECC_REG_ECC_MSG_1                                                                       (32'h10008104)
`define ECC_REG_ECC_MSG_1                                                                           (32'h104)
`define CLP_ECC_REG_ECC_MSG_2                                                                       (32'h10008108)
`define ECC_REG_ECC_MSG_2                                                                           (32'h108)
`define CLP_ECC_REG_ECC_MSG_3                                                                       (32'h1000810c)
`define ECC_REG_ECC_MSG_3                                                                           (32'h10c)
`define CLP_ECC_REG_ECC_MSG_4                                                                       (32'h10008110)
`define ECC_REG_ECC_MSG_4                                                                           (32'h110)
`define CLP_ECC_REG_ECC_MSG_5                                                                       (32'h10008114)
`define ECC_REG_ECC_MSG_5                                                                           (32'h114)
`define CLP_ECC_REG_ECC_MSG_6                                                                       (32'h10008118)
`define ECC_REG_ECC_MSG_6                                                                           (32'h118)
`define CLP_ECC_REG_ECC_MSG_7                                                                       (32'h1000811c)
`define ECC_REG_ECC_MSG_7                                                                           (32'h11c)
`define CLP_ECC_REG_ECC_MSG_8                                                                       (32'h10008120)
`define ECC_REG_ECC_MSG_8                                                                           (32'h120)
`define CLP_ECC_REG_ECC_MSG_9                                                                       (32'h10008124)
`define ECC_REG_ECC_MSG_9                                                                           (32'h124)
`define CLP_ECC_REG_ECC_MSG_10                                                                      (32'h10008128)
`define ECC_REG_ECC_MSG_10                                                                          (32'h128)
`define CLP_ECC_REG_ECC_MSG_11                                                                      (32'h1000812c)
`define ECC_REG_ECC_MSG_11                                                                          (32'h12c)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_0                                                               (32'h10008180)
`define ECC_REG_ECC_PRIVKEY_OUT_0                                                                   (32'h180)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_1                                                               (32'h10008184)
`define ECC_REG_ECC_PRIVKEY_OUT_1                                                                   (32'h184)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_2                                                               (32'h10008188)
`define ECC_REG_ECC_PRIVKEY_OUT_2                                                                   (32'h188)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_3                                                               (32'h1000818c)
`define ECC_REG_ECC_PRIVKEY_OUT_3                                                                   (32'h18c)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_4                                                               (32'h10008190)
`define ECC_REG_ECC_PRIVKEY_OUT_4                                                                   (32'h190)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_5                                                               (32'h10008194)
`define ECC_REG_ECC_PRIVKEY_OUT_5                                                                   (32'h194)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_6                                                               (32'h10008198)
`define ECC_REG_ECC_PRIVKEY_OUT_6                                                                   (32'h198)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_7                                                               (32'h1000819c)
`define ECC_REG_ECC_PRIVKEY_OUT_7                                                                   (32'h19c)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_8                                                               (32'h100081a0)
`define ECC_REG_ECC_PRIVKEY_OUT_8                                                                   (32'h1a0)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_9                                                               (32'h100081a4)
`define ECC_REG_ECC_PRIVKEY_OUT_9                                                                   (32'h1a4)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_10                                                              (32'h100081a8)
`define ECC_REG_ECC_PRIVKEY_OUT_10                                                                  (32'h1a8)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_11                                                              (32'h100081ac)
`define ECC_REG_ECC_PRIVKEY_OUT_11                                                                  (32'h1ac)
`define CLP_ECC_REG_ECC_PUBKEY_X_0                                                                  (32'h10008200)
`define ECC_REG_ECC_PUBKEY_X_0                                                                      (32'h200)
`define CLP_ECC_REG_ECC_PUBKEY_X_1                                                                  (32'h10008204)
`define ECC_REG_ECC_PUBKEY_X_1                                                                      (32'h204)
`define CLP_ECC_REG_ECC_PUBKEY_X_2                                                                  (32'h10008208)
`define ECC_REG_ECC_PUBKEY_X_2                                                                      (32'h208)
`define CLP_ECC_REG_ECC_PUBKEY_X_3                                                                  (32'h1000820c)
`define ECC_REG_ECC_PUBKEY_X_3                                                                      (32'h20c)
`define CLP_ECC_REG_ECC_PUBKEY_X_4                                                                  (32'h10008210)
`define ECC_REG_ECC_PUBKEY_X_4                                                                      (32'h210)
`define CLP_ECC_REG_ECC_PUBKEY_X_5                                                                  (32'h10008214)
`define ECC_REG_ECC_PUBKEY_X_5                                                                      (32'h214)
`define CLP_ECC_REG_ECC_PUBKEY_X_6                                                                  (32'h10008218)
`define ECC_REG_ECC_PUBKEY_X_6                                                                      (32'h218)
`define CLP_ECC_REG_ECC_PUBKEY_X_7                                                                  (32'h1000821c)
`define ECC_REG_ECC_PUBKEY_X_7                                                                      (32'h21c)
`define CLP_ECC_REG_ECC_PUBKEY_X_8                                                                  (32'h10008220)
`define ECC_REG_ECC_PUBKEY_X_8                                                                      (32'h220)
`define CLP_ECC_REG_ECC_PUBKEY_X_9                                                                  (32'h10008224)
`define ECC_REG_ECC_PUBKEY_X_9                                                                      (32'h224)
`define CLP_ECC_REG_ECC_PUBKEY_X_10                                                                 (32'h10008228)
`define ECC_REG_ECC_PUBKEY_X_10                                                                     (32'h228)
`define CLP_ECC_REG_ECC_PUBKEY_X_11                                                                 (32'h1000822c)
`define ECC_REG_ECC_PUBKEY_X_11                                                                     (32'h22c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_0                                                                  (32'h10008280)
`define ECC_REG_ECC_PUBKEY_Y_0                                                                      (32'h280)
`define CLP_ECC_REG_ECC_PUBKEY_Y_1                                                                  (32'h10008284)
`define ECC_REG_ECC_PUBKEY_Y_1                                                                      (32'h284)
`define CLP_ECC_REG_ECC_PUBKEY_Y_2                                                                  (32'h10008288)
`define ECC_REG_ECC_PUBKEY_Y_2                                                                      (32'h288)
`define CLP_ECC_REG_ECC_PUBKEY_Y_3                                                                  (32'h1000828c)
`define ECC_REG_ECC_PUBKEY_Y_3                                                                      (32'h28c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_4                                                                  (32'h10008290)
`define ECC_REG_ECC_PUBKEY_Y_4                                                                      (32'h290)
`define CLP_ECC_REG_ECC_PUBKEY_Y_5                                                                  (32'h10008294)
`define ECC_REG_ECC_PUBKEY_Y_5                                                                      (32'h294)
`define CLP_ECC_REG_ECC_PUBKEY_Y_6                                                                  (32'h10008298)
`define ECC_REG_ECC_PUBKEY_Y_6                                                                      (32'h298)
`define CLP_ECC_REG_ECC_PUBKEY_Y_7                                                                  (32'h1000829c)
`define ECC_REG_ECC_PUBKEY_Y_7                                                                      (32'h29c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_8                                                                  (32'h100082a0)
`define ECC_REG_ECC_PUBKEY_Y_8                                                                      (32'h2a0)
`define CLP_ECC_REG_ECC_PUBKEY_Y_9                                                                  (32'h100082a4)
`define ECC_REG_ECC_PUBKEY_Y_9                                                                      (32'h2a4)
`define CLP_ECC_REG_ECC_PUBKEY_Y_10                                                                 (32'h100082a8)
`define ECC_REG_ECC_PUBKEY_Y_10                                                                     (32'h2a8)
`define CLP_ECC_REG_ECC_PUBKEY_Y_11                                                                 (32'h100082ac)
`define ECC_REG_ECC_PUBKEY_Y_11                                                                     (32'h2ac)
`define CLP_ECC_REG_ECC_SIGN_R_0                                                                    (32'h10008300)
`define ECC_REG_ECC_SIGN_R_0                                                                        (32'h300)
`define CLP_ECC_REG_ECC_SIGN_R_1                                                                    (32'h10008304)
`define ECC_REG_ECC_SIGN_R_1                                                                        (32'h304)
`define CLP_ECC_REG_ECC_SIGN_R_2                                                                    (32'h10008308)
`define ECC_REG_ECC_SIGN_R_2                                                                        (32'h308)
`define CLP_ECC_REG_ECC_SIGN_R_3                                                                    (32'h1000830c)
`define ECC_REG_ECC_SIGN_R_3                                                                        (32'h30c)
`define CLP_ECC_REG_ECC_SIGN_R_4                                                                    (32'h10008310)
`define ECC_REG_ECC_SIGN_R_4                                                                        (32'h310)
`define CLP_ECC_REG_ECC_SIGN_R_5                                                                    (32'h10008314)
`define ECC_REG_ECC_SIGN_R_5                                                                        (32'h314)
`define CLP_ECC_REG_ECC_SIGN_R_6                                                                    (32'h10008318)
`define ECC_REG_ECC_SIGN_R_6                                                                        (32'h318)
`define CLP_ECC_REG_ECC_SIGN_R_7                                                                    (32'h1000831c)
`define ECC_REG_ECC_SIGN_R_7                                                                        (32'h31c)
`define CLP_ECC_REG_ECC_SIGN_R_8                                                                    (32'h10008320)
`define ECC_REG_ECC_SIGN_R_8                                                                        (32'h320)
`define CLP_ECC_REG_ECC_SIGN_R_9                                                                    (32'h10008324)
`define ECC_REG_ECC_SIGN_R_9                                                                        (32'h324)
`define CLP_ECC_REG_ECC_SIGN_R_10                                                                   (32'h10008328)
`define ECC_REG_ECC_SIGN_R_10                                                                       (32'h328)
`define CLP_ECC_REG_ECC_SIGN_R_11                                                                   (32'h1000832c)
`define ECC_REG_ECC_SIGN_R_11                                                                       (32'h32c)
`define CLP_ECC_REG_ECC_SIGN_S_0                                                                    (32'h10008380)
`define ECC_REG_ECC_SIGN_S_0                                                                        (32'h380)
`define CLP_ECC_REG_ECC_SIGN_S_1                                                                    (32'h10008384)
`define ECC_REG_ECC_SIGN_S_1                                                                        (32'h384)
`define CLP_ECC_REG_ECC_SIGN_S_2                                                                    (32'h10008388)
`define ECC_REG_ECC_SIGN_S_2                                                                        (32'h388)
`define CLP_ECC_REG_ECC_SIGN_S_3                                                                    (32'h1000838c)
`define ECC_REG_ECC_SIGN_S_3                                                                        (32'h38c)
`define CLP_ECC_REG_ECC_SIGN_S_4                                                                    (32'h10008390)
`define ECC_REG_ECC_SIGN_S_4                                                                        (32'h390)
`define CLP_ECC_REG_ECC_SIGN_S_5                                                                    (32'h10008394)
`define ECC_REG_ECC_SIGN_S_5                                                                        (32'h394)
`define CLP_ECC_REG_ECC_SIGN_S_6                                                                    (32'h10008398)
`define ECC_REG_ECC_SIGN_S_6                                                                        (32'h398)
`define CLP_ECC_REG_ECC_SIGN_S_7                                                                    (32'h1000839c)
`define ECC_REG_ECC_SIGN_S_7                                                                        (32'h39c)
`define CLP_ECC_REG_ECC_SIGN_S_8                                                                    (32'h100083a0)
`define ECC_REG_ECC_SIGN_S_8                                                                        (32'h3a0)
`define CLP_ECC_REG_ECC_SIGN_S_9                                                                    (32'h100083a4)
`define ECC_REG_ECC_SIGN_S_9                                                                        (32'h3a4)
`define CLP_ECC_REG_ECC_SIGN_S_10                                                                   (32'h100083a8)
`define ECC_REG_ECC_SIGN_S_10                                                                       (32'h3a8)
`define CLP_ECC_REG_ECC_SIGN_S_11                                                                   (32'h100083ac)
`define ECC_REG_ECC_SIGN_S_11                                                                       (32'h3ac)
`define CLP_ECC_REG_ECC_VERIFY_R_0                                                                  (32'h10008400)
`define ECC_REG_ECC_VERIFY_R_0                                                                      (32'h400)
`define CLP_ECC_REG_ECC_VERIFY_R_1                                                                  (32'h10008404)
`define ECC_REG_ECC_VERIFY_R_1                                                                      (32'h404)
`define CLP_ECC_REG_ECC_VERIFY_R_2                                                                  (32'h10008408)
`define ECC_REG_ECC_VERIFY_R_2                                                                      (32'h408)
`define CLP_ECC_REG_ECC_VERIFY_R_3                                                                  (32'h1000840c)
`define ECC_REG_ECC_VERIFY_R_3                                                                      (32'h40c)
`define CLP_ECC_REG_ECC_VERIFY_R_4                                                                  (32'h10008410)
`define ECC_REG_ECC_VERIFY_R_4                                                                      (32'h410)
`define CLP_ECC_REG_ECC_VERIFY_R_5                                                                  (32'h10008414)
`define ECC_REG_ECC_VERIFY_R_5                                                                      (32'h414)
`define CLP_ECC_REG_ECC_VERIFY_R_6                                                                  (32'h10008418)
`define ECC_REG_ECC_VERIFY_R_6                                                                      (32'h418)
`define CLP_ECC_REG_ECC_VERIFY_R_7                                                                  (32'h1000841c)
`define ECC_REG_ECC_VERIFY_R_7                                                                      (32'h41c)
`define CLP_ECC_REG_ECC_VERIFY_R_8                                                                  (32'h10008420)
`define ECC_REG_ECC_VERIFY_R_8                                                                      (32'h420)
`define CLP_ECC_REG_ECC_VERIFY_R_9                                                                  (32'h10008424)
`define ECC_REG_ECC_VERIFY_R_9                                                                      (32'h424)
`define CLP_ECC_REG_ECC_VERIFY_R_10                                                                 (32'h10008428)
`define ECC_REG_ECC_VERIFY_R_10                                                                     (32'h428)
`define CLP_ECC_REG_ECC_VERIFY_R_11                                                                 (32'h1000842c)
`define ECC_REG_ECC_VERIFY_R_11                                                                     (32'h42c)
`define CLP_ECC_REG_ECC_IV_0                                                                        (32'h10008480)
`define ECC_REG_ECC_IV_0                                                                            (32'h480)
`define CLP_ECC_REG_ECC_IV_1                                                                        (32'h10008484)
`define ECC_REG_ECC_IV_1                                                                            (32'h484)
`define CLP_ECC_REG_ECC_IV_2                                                                        (32'h10008488)
`define ECC_REG_ECC_IV_2                                                                            (32'h488)
`define CLP_ECC_REG_ECC_IV_3                                                                        (32'h1000848c)
`define ECC_REG_ECC_IV_3                                                                            (32'h48c)
`define CLP_ECC_REG_ECC_IV_4                                                                        (32'h10008490)
`define ECC_REG_ECC_IV_4                                                                            (32'h490)
`define CLP_ECC_REG_ECC_IV_5                                                                        (32'h10008494)
`define ECC_REG_ECC_IV_5                                                                            (32'h494)
`define CLP_ECC_REG_ECC_IV_6                                                                        (32'h10008498)
`define ECC_REG_ECC_IV_6                                                                            (32'h498)
`define CLP_ECC_REG_ECC_IV_7                                                                        (32'h1000849c)
`define ECC_REG_ECC_IV_7                                                                            (32'h49c)
`define CLP_ECC_REG_ECC_IV_8                                                                        (32'h100084a0)
`define ECC_REG_ECC_IV_8                                                                            (32'h4a0)
`define CLP_ECC_REG_ECC_IV_9                                                                        (32'h100084a4)
`define ECC_REG_ECC_IV_9                                                                            (32'h4a4)
`define CLP_ECC_REG_ECC_IV_10                                                                       (32'h100084a8)
`define ECC_REG_ECC_IV_10                                                                           (32'h4a8)
`define CLP_ECC_REG_ECC_IV_11                                                                       (32'h100084ac)
`define ECC_REG_ECC_IV_11                                                                           (32'h4ac)
`define CLP_ECC_REG_ECC_NONCE_0                                                                     (32'h10008500)
`define ECC_REG_ECC_NONCE_0                                                                         (32'h500)
`define CLP_ECC_REG_ECC_NONCE_1                                                                     (32'h10008504)
`define ECC_REG_ECC_NONCE_1                                                                         (32'h504)
`define CLP_ECC_REG_ECC_NONCE_2                                                                     (32'h10008508)
`define ECC_REG_ECC_NONCE_2                                                                         (32'h508)
`define CLP_ECC_REG_ECC_NONCE_3                                                                     (32'h1000850c)
`define ECC_REG_ECC_NONCE_3                                                                         (32'h50c)
`define CLP_ECC_REG_ECC_NONCE_4                                                                     (32'h10008510)
`define ECC_REG_ECC_NONCE_4                                                                         (32'h510)
`define CLP_ECC_REG_ECC_NONCE_5                                                                     (32'h10008514)
`define ECC_REG_ECC_NONCE_5                                                                         (32'h514)
`define CLP_ECC_REG_ECC_NONCE_6                                                                     (32'h10008518)
`define ECC_REG_ECC_NONCE_6                                                                         (32'h518)
`define CLP_ECC_REG_ECC_NONCE_7                                                                     (32'h1000851c)
`define ECC_REG_ECC_NONCE_7                                                                         (32'h51c)
`define CLP_ECC_REG_ECC_NONCE_8                                                                     (32'h10008520)
`define ECC_REG_ECC_NONCE_8                                                                         (32'h520)
`define CLP_ECC_REG_ECC_NONCE_9                                                                     (32'h10008524)
`define ECC_REG_ECC_NONCE_9                                                                         (32'h524)
`define CLP_ECC_REG_ECC_NONCE_10                                                                    (32'h10008528)
`define ECC_REG_ECC_NONCE_10                                                                        (32'h528)
`define CLP_ECC_REG_ECC_NONCE_11                                                                    (32'h1000852c)
`define ECC_REG_ECC_NONCE_11                                                                        (32'h52c)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_0                                                                (32'h10008580)
`define ECC_REG_ECC_PRIVKEY_IN_0                                                                    (32'h580)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_1                                                                (32'h10008584)
`define ECC_REG_ECC_PRIVKEY_IN_1                                                                    (32'h584)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_2                                                                (32'h10008588)
`define ECC_REG_ECC_PRIVKEY_IN_2                                                                    (32'h588)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_3                                                                (32'h1000858c)
`define ECC_REG_ECC_PRIVKEY_IN_3                                                                    (32'h58c)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_4                                                                (32'h10008590)
`define ECC_REG_ECC_PRIVKEY_IN_4                                                                    (32'h590)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_5                                                                (32'h10008594)
`define ECC_REG_ECC_PRIVKEY_IN_5                                                                    (32'h594)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_6                                                                (32'h10008598)
`define ECC_REG_ECC_PRIVKEY_IN_6                                                                    (32'h598)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_7                                                                (32'h1000859c)
`define ECC_REG_ECC_PRIVKEY_IN_7                                                                    (32'h59c)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_8                                                                (32'h100085a0)
`define ECC_REG_ECC_PRIVKEY_IN_8                                                                    (32'h5a0)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_9                                                                (32'h100085a4)
`define ECC_REG_ECC_PRIVKEY_IN_9                                                                    (32'h5a4)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_10                                                               (32'h100085a8)
`define ECC_REG_ECC_PRIVKEY_IN_10                                                                   (32'h5a8)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_11                                                               (32'h100085ac)
`define ECC_REG_ECC_PRIVKEY_IN_11                                                                   (32'h5ac)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_0                                                             (32'h100085c0)
`define ECC_REG_ECC_DH_SHARED_KEY_0                                                                 (32'h5c0)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_1                                                             (32'h100085c4)
`define ECC_REG_ECC_DH_SHARED_KEY_1                                                                 (32'h5c4)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_2                                                             (32'h100085c8)
`define ECC_REG_ECC_DH_SHARED_KEY_2                                                                 (32'h5c8)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_3                                                             (32'h100085cc)
`define ECC_REG_ECC_DH_SHARED_KEY_3                                                                 (32'h5cc)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_4                                                             (32'h100085d0)
`define ECC_REG_ECC_DH_SHARED_KEY_4                                                                 (32'h5d0)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_5                                                             (32'h100085d4)
`define ECC_REG_ECC_DH_SHARED_KEY_5                                                                 (32'h5d4)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_6                                                             (32'h100085d8)
`define ECC_REG_ECC_DH_SHARED_KEY_6                                                                 (32'h5d8)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_7                                                             (32'h100085dc)
`define ECC_REG_ECC_DH_SHARED_KEY_7                                                                 (32'h5dc)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_8                                                             (32'h100085e0)
`define ECC_REG_ECC_DH_SHARED_KEY_8                                                                 (32'h5e0)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_9                                                             (32'h100085e4)
`define ECC_REG_ECC_DH_SHARED_KEY_9                                                                 (32'h5e4)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_10                                                            (32'h100085e8)
`define ECC_REG_ECC_DH_SHARED_KEY_10                                                                (32'h5e8)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_11                                                            (32'h100085ec)
`define ECC_REG_ECC_DH_SHARED_KEY_11                                                                (32'h5ec)
`define CLP_ECC_REG_ECC_KV_RD_PKEY_CTRL                                                             (32'h10008600)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL                                                                 (32'h600)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_EN_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_EN_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_ENTRY_LOW                                                  (1)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_ENTRY_MASK                                                 (32'h3e)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_PCR_HASH_EXTEND_LOW                                             (6)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_PCR_HASH_EXTEND_MASK                                            (32'h40)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_RSVD_LOW                                                        (7)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_RSVD_MASK                                                       (32'hffffff80)
`define CLP_ECC_REG_ECC_KV_RD_PKEY_STATUS                                                           (32'h10008604)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS                                                               (32'h604)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_ECC_KV_RD_SEED_CTRL                                                             (32'h10008608)
`define ECC_REG_ECC_KV_RD_SEED_CTRL                                                                 (32'h608)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_EN_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_EN_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_ENTRY_LOW                                                  (1)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_ENTRY_MASK                                                 (32'h3e)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_PCR_HASH_EXTEND_LOW                                             (6)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_PCR_HASH_EXTEND_MASK                                            (32'h40)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_RSVD_LOW                                                        (7)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_RSVD_MASK                                                       (32'hffffff80)
`define CLP_ECC_REG_ECC_KV_RD_SEED_STATUS                                                           (32'h1000860c)
`define ECC_REG_ECC_KV_RD_SEED_STATUS                                                               (32'h60c)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_ECC_KV_WR_PKEY_CTRL                                                             (32'h10008610)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL                                                                 (32'h610)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_EN_LOW                                                    (0)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_EN_MASK                                                   (32'h1)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_ENTRY_LOW                                                 (1)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_ENTRY_MASK                                                (32'h3e)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_KEY_DEST_VALID_LOW                                         (6)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_KEY_DEST_VALID_MASK                                        (32'h40)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                       (7)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                      (32'h80)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_SHA_BLOCK_DEST_VALID_LOW                                        (8)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_SHA_BLOCK_DEST_VALID_MASK                                       (32'h100)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_PKEY_DEST_VALID_LOW                                         (9)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_PKEY_DEST_VALID_MASK                                        (32'h200)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_SEED_DEST_VALID_LOW                                         (10)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_SEED_DEST_VALID_MASK                                        (32'h400)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_RSVD_LOW                                                        (11)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_RSVD_MASK                                                       (32'hfffff800)
`define CLP_ECC_REG_ECC_KV_WR_PKEY_STATUS                                                           (32'h10008614)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS                                                               (32'h614)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_INTR_BLOCK_RF_START                                                             (32'h10008800)
`define CLP_ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10008800)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                      (32'h800)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                         (0)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                        (32'h1)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                         (1)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                        (32'h2)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10008804)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                       (32'h804)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_LOW                                 (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_MASK                                (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10008808)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                       (32'h808)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                 (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                                (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1000880c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                   (32'h80c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10008810)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                   (32'h810)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10008814)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                 (32'h814)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_LOW                          (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_MASK                         (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10008818)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                 (32'h818)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                          (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                         (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1000881c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                     (32'h81c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_LOW                             (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_MASK                            (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10008820)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                     (32'h820)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                             (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                            (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h10008900)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                           (32'h900)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10008980)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                           (32'h980)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'h10008a00)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                      (32'ha00)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10008a04)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                      (32'ha04)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_HMAC_REG_BASE_ADDR                                                                      (32'h10010000)
`define CLP_HMAC_REG_HMAC512_NAME_0                                                                 (32'h10010000)
`define HMAC_REG_HMAC512_NAME_0                                                                     (32'h0)
`define CLP_HMAC_REG_HMAC512_NAME_1                                                                 (32'h10010004)
`define HMAC_REG_HMAC512_NAME_1                                                                     (32'h4)
`define CLP_HMAC_REG_HMAC512_VERSION_0                                                              (32'h10010008)
`define HMAC_REG_HMAC512_VERSION_0                                                                  (32'h8)
`define CLP_HMAC_REG_HMAC512_VERSION_1                                                              (32'h1001000c)
`define HMAC_REG_HMAC512_VERSION_1                                                                  (32'hc)
`define CLP_HMAC_REG_HMAC512_CTRL                                                                   (32'h10010010)
`define HMAC_REG_HMAC512_CTRL                                                                       (32'h10)
`define HMAC_REG_HMAC512_CTRL_INIT_LOW                                                              (0)
`define HMAC_REG_HMAC512_CTRL_INIT_MASK                                                             (32'h1)
`define HMAC_REG_HMAC512_CTRL_NEXT_LOW                                                              (1)
`define HMAC_REG_HMAC512_CTRL_NEXT_MASK                                                             (32'h2)
`define HMAC_REG_HMAC512_CTRL_ZEROIZE_LOW                                                           (2)
`define HMAC_REG_HMAC512_CTRL_ZEROIZE_MASK                                                          (32'h4)
`define HMAC_REG_HMAC512_CTRL_MODE_LOW                                                              (3)
`define HMAC_REG_HMAC512_CTRL_MODE_MASK                                                             (32'h8)
`define HMAC_REG_HMAC512_CTRL_RESERVED_LOW                                                          (4)
`define HMAC_REG_HMAC512_CTRL_RESERVED_MASK                                                         (32'h10)
`define CLP_HMAC_REG_HMAC512_STATUS                                                                 (32'h10010018)
`define HMAC_REG_HMAC512_STATUS                                                                     (32'h18)
`define HMAC_REG_HMAC512_STATUS_READY_LOW                                                           (0)
`define HMAC_REG_HMAC512_STATUS_READY_MASK                                                          (32'h1)
`define HMAC_REG_HMAC512_STATUS_VALID_LOW                                                           (1)
`define HMAC_REG_HMAC512_STATUS_VALID_MASK                                                          (32'h2)
`define CLP_HMAC_REG_HMAC512_KEY_0                                                                  (32'h10010040)
`define HMAC_REG_HMAC512_KEY_0                                                                      (32'h40)
`define CLP_HMAC_REG_HMAC512_KEY_1                                                                  (32'h10010044)
`define HMAC_REG_HMAC512_KEY_1                                                                      (32'h44)
`define CLP_HMAC_REG_HMAC512_KEY_2                                                                  (32'h10010048)
`define HMAC_REG_HMAC512_KEY_2                                                                      (32'h48)
`define CLP_HMAC_REG_HMAC512_KEY_3                                                                  (32'h1001004c)
`define HMAC_REG_HMAC512_KEY_3                                                                      (32'h4c)
`define CLP_HMAC_REG_HMAC512_KEY_4                                                                  (32'h10010050)
`define HMAC_REG_HMAC512_KEY_4                                                                      (32'h50)
`define CLP_HMAC_REG_HMAC512_KEY_5                                                                  (32'h10010054)
`define HMAC_REG_HMAC512_KEY_5                                                                      (32'h54)
`define CLP_HMAC_REG_HMAC512_KEY_6                                                                  (32'h10010058)
`define HMAC_REG_HMAC512_KEY_6                                                                      (32'h58)
`define CLP_HMAC_REG_HMAC512_KEY_7                                                                  (32'h1001005c)
`define HMAC_REG_HMAC512_KEY_7                                                                      (32'h5c)
`define CLP_HMAC_REG_HMAC512_KEY_8                                                                  (32'h10010060)
`define HMAC_REG_HMAC512_KEY_8                                                                      (32'h60)
`define CLP_HMAC_REG_HMAC512_KEY_9                                                                  (32'h10010064)
`define HMAC_REG_HMAC512_KEY_9                                                                      (32'h64)
`define CLP_HMAC_REG_HMAC512_KEY_10                                                                 (32'h10010068)
`define HMAC_REG_HMAC512_KEY_10                                                                     (32'h68)
`define CLP_HMAC_REG_HMAC512_KEY_11                                                                 (32'h1001006c)
`define HMAC_REG_HMAC512_KEY_11                                                                     (32'h6c)
`define CLP_HMAC_REG_HMAC512_KEY_12                                                                 (32'h10010070)
`define HMAC_REG_HMAC512_KEY_12                                                                     (32'h70)
`define CLP_HMAC_REG_HMAC512_KEY_13                                                                 (32'h10010074)
`define HMAC_REG_HMAC512_KEY_13                                                                     (32'h74)
`define CLP_HMAC_REG_HMAC512_KEY_14                                                                 (32'h10010078)
`define HMAC_REG_HMAC512_KEY_14                                                                     (32'h78)
`define CLP_HMAC_REG_HMAC512_KEY_15                                                                 (32'h1001007c)
`define HMAC_REG_HMAC512_KEY_15                                                                     (32'h7c)
`define CLP_HMAC_REG_HMAC512_BLOCK_0                                                                (32'h10010080)
`define HMAC_REG_HMAC512_BLOCK_0                                                                    (32'h80)
`define CLP_HMAC_REG_HMAC512_BLOCK_1                                                                (32'h10010084)
`define HMAC_REG_HMAC512_BLOCK_1                                                                    (32'h84)
`define CLP_HMAC_REG_HMAC512_BLOCK_2                                                                (32'h10010088)
`define HMAC_REG_HMAC512_BLOCK_2                                                                    (32'h88)
`define CLP_HMAC_REG_HMAC512_BLOCK_3                                                                (32'h1001008c)
`define HMAC_REG_HMAC512_BLOCK_3                                                                    (32'h8c)
`define CLP_HMAC_REG_HMAC512_BLOCK_4                                                                (32'h10010090)
`define HMAC_REG_HMAC512_BLOCK_4                                                                    (32'h90)
`define CLP_HMAC_REG_HMAC512_BLOCK_5                                                                (32'h10010094)
`define HMAC_REG_HMAC512_BLOCK_5                                                                    (32'h94)
`define CLP_HMAC_REG_HMAC512_BLOCK_6                                                                (32'h10010098)
`define HMAC_REG_HMAC512_BLOCK_6                                                                    (32'h98)
`define CLP_HMAC_REG_HMAC512_BLOCK_7                                                                (32'h1001009c)
`define HMAC_REG_HMAC512_BLOCK_7                                                                    (32'h9c)
`define CLP_HMAC_REG_HMAC512_BLOCK_8                                                                (32'h100100a0)
`define HMAC_REG_HMAC512_BLOCK_8                                                                    (32'ha0)
`define CLP_HMAC_REG_HMAC512_BLOCK_9                                                                (32'h100100a4)
`define HMAC_REG_HMAC512_BLOCK_9                                                                    (32'ha4)
`define CLP_HMAC_REG_HMAC512_BLOCK_10                                                               (32'h100100a8)
`define HMAC_REG_HMAC512_BLOCK_10                                                                   (32'ha8)
`define CLP_HMAC_REG_HMAC512_BLOCK_11                                                               (32'h100100ac)
`define HMAC_REG_HMAC512_BLOCK_11                                                                   (32'hac)
`define CLP_HMAC_REG_HMAC512_BLOCK_12                                                               (32'h100100b0)
`define HMAC_REG_HMAC512_BLOCK_12                                                                   (32'hb0)
`define CLP_HMAC_REG_HMAC512_BLOCK_13                                                               (32'h100100b4)
`define HMAC_REG_HMAC512_BLOCK_13                                                                   (32'hb4)
`define CLP_HMAC_REG_HMAC512_BLOCK_14                                                               (32'h100100b8)
`define HMAC_REG_HMAC512_BLOCK_14                                                                   (32'hb8)
`define CLP_HMAC_REG_HMAC512_BLOCK_15                                                               (32'h100100bc)
`define HMAC_REG_HMAC512_BLOCK_15                                                                   (32'hbc)
`define CLP_HMAC_REG_HMAC512_BLOCK_16                                                               (32'h100100c0)
`define HMAC_REG_HMAC512_BLOCK_16                                                                   (32'hc0)
`define CLP_HMAC_REG_HMAC512_BLOCK_17                                                               (32'h100100c4)
`define HMAC_REG_HMAC512_BLOCK_17                                                                   (32'hc4)
`define CLP_HMAC_REG_HMAC512_BLOCK_18                                                               (32'h100100c8)
`define HMAC_REG_HMAC512_BLOCK_18                                                                   (32'hc8)
`define CLP_HMAC_REG_HMAC512_BLOCK_19                                                               (32'h100100cc)
`define HMAC_REG_HMAC512_BLOCK_19                                                                   (32'hcc)
`define CLP_HMAC_REG_HMAC512_BLOCK_20                                                               (32'h100100d0)
`define HMAC_REG_HMAC512_BLOCK_20                                                                   (32'hd0)
`define CLP_HMAC_REG_HMAC512_BLOCK_21                                                               (32'h100100d4)
`define HMAC_REG_HMAC512_BLOCK_21                                                                   (32'hd4)
`define CLP_HMAC_REG_HMAC512_BLOCK_22                                                               (32'h100100d8)
`define HMAC_REG_HMAC512_BLOCK_22                                                                   (32'hd8)
`define CLP_HMAC_REG_HMAC512_BLOCK_23                                                               (32'h100100dc)
`define HMAC_REG_HMAC512_BLOCK_23                                                                   (32'hdc)
`define CLP_HMAC_REG_HMAC512_BLOCK_24                                                               (32'h100100e0)
`define HMAC_REG_HMAC512_BLOCK_24                                                                   (32'he0)
`define CLP_HMAC_REG_HMAC512_BLOCK_25                                                               (32'h100100e4)
`define HMAC_REG_HMAC512_BLOCK_25                                                                   (32'he4)
`define CLP_HMAC_REG_HMAC512_BLOCK_26                                                               (32'h100100e8)
`define HMAC_REG_HMAC512_BLOCK_26                                                                   (32'he8)
`define CLP_HMAC_REG_HMAC512_BLOCK_27                                                               (32'h100100ec)
`define HMAC_REG_HMAC512_BLOCK_27                                                                   (32'hec)
`define CLP_HMAC_REG_HMAC512_BLOCK_28                                                               (32'h100100f0)
`define HMAC_REG_HMAC512_BLOCK_28                                                                   (32'hf0)
`define CLP_HMAC_REG_HMAC512_BLOCK_29                                                               (32'h100100f4)
`define HMAC_REG_HMAC512_BLOCK_29                                                                   (32'hf4)
`define CLP_HMAC_REG_HMAC512_BLOCK_30                                                               (32'h100100f8)
`define HMAC_REG_HMAC512_BLOCK_30                                                                   (32'hf8)
`define CLP_HMAC_REG_HMAC512_BLOCK_31                                                               (32'h100100fc)
`define HMAC_REG_HMAC512_BLOCK_31                                                                   (32'hfc)
`define CLP_HMAC_REG_HMAC512_TAG_0                                                                  (32'h10010100)
`define HMAC_REG_HMAC512_TAG_0                                                                      (32'h100)
`define CLP_HMAC_REG_HMAC512_TAG_1                                                                  (32'h10010104)
`define HMAC_REG_HMAC512_TAG_1                                                                      (32'h104)
`define CLP_HMAC_REG_HMAC512_TAG_2                                                                  (32'h10010108)
`define HMAC_REG_HMAC512_TAG_2                                                                      (32'h108)
`define CLP_HMAC_REG_HMAC512_TAG_3                                                                  (32'h1001010c)
`define HMAC_REG_HMAC512_TAG_3                                                                      (32'h10c)
`define CLP_HMAC_REG_HMAC512_TAG_4                                                                  (32'h10010110)
`define HMAC_REG_HMAC512_TAG_4                                                                      (32'h110)
`define CLP_HMAC_REG_HMAC512_TAG_5                                                                  (32'h10010114)
`define HMAC_REG_HMAC512_TAG_5                                                                      (32'h114)
`define CLP_HMAC_REG_HMAC512_TAG_6                                                                  (32'h10010118)
`define HMAC_REG_HMAC512_TAG_6                                                                      (32'h118)
`define CLP_HMAC_REG_HMAC512_TAG_7                                                                  (32'h1001011c)
`define HMAC_REG_HMAC512_TAG_7                                                                      (32'h11c)
`define CLP_HMAC_REG_HMAC512_TAG_8                                                                  (32'h10010120)
`define HMAC_REG_HMAC512_TAG_8                                                                      (32'h120)
`define CLP_HMAC_REG_HMAC512_TAG_9                                                                  (32'h10010124)
`define HMAC_REG_HMAC512_TAG_9                                                                      (32'h124)
`define CLP_HMAC_REG_HMAC512_TAG_10                                                                 (32'h10010128)
`define HMAC_REG_HMAC512_TAG_10                                                                     (32'h128)
`define CLP_HMAC_REG_HMAC512_TAG_11                                                                 (32'h1001012c)
`define HMAC_REG_HMAC512_TAG_11                                                                     (32'h12c)
`define CLP_HMAC_REG_HMAC512_TAG_12                                                                 (32'h10010130)
`define HMAC_REG_HMAC512_TAG_12                                                                     (32'h130)
`define CLP_HMAC_REG_HMAC512_TAG_13                                                                 (32'h10010134)
`define HMAC_REG_HMAC512_TAG_13                                                                     (32'h134)
`define CLP_HMAC_REG_HMAC512_TAG_14                                                                 (32'h10010138)
`define HMAC_REG_HMAC512_TAG_14                                                                     (32'h138)
`define CLP_HMAC_REG_HMAC512_TAG_15                                                                 (32'h1001013c)
`define HMAC_REG_HMAC512_TAG_15                                                                     (32'h13c)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_0                                                            (32'h10010130)
`define HMAC_REG_HMAC512_LFSR_SEED_0                                                                (32'h130)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_1                                                            (32'h10010134)
`define HMAC_REG_HMAC512_LFSR_SEED_1                                                                (32'h134)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_2                                                            (32'h10010138)
`define HMAC_REG_HMAC512_LFSR_SEED_2                                                                (32'h138)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_3                                                            (32'h1001013c)
`define HMAC_REG_HMAC512_LFSR_SEED_3                                                                (32'h13c)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_4                                                            (32'h10010140)
`define HMAC_REG_HMAC512_LFSR_SEED_4                                                                (32'h140)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_5                                                            (32'h10010144)
`define HMAC_REG_HMAC512_LFSR_SEED_5                                                                (32'h144)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_6                                                            (32'h10010148)
`define HMAC_REG_HMAC512_LFSR_SEED_6                                                                (32'h148)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_7                                                            (32'h1001014c)
`define HMAC_REG_HMAC512_LFSR_SEED_7                                                                (32'h14c)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_8                                                            (32'h10010150)
`define HMAC_REG_HMAC512_LFSR_SEED_8                                                                (32'h150)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_9                                                            (32'h10010154)
`define HMAC_REG_HMAC512_LFSR_SEED_9                                                                (32'h154)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_10                                                           (32'h10010158)
`define HMAC_REG_HMAC512_LFSR_SEED_10                                                               (32'h158)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_11                                                           (32'h1001015c)
`define HMAC_REG_HMAC512_LFSR_SEED_11                                                               (32'h15c)
`define CLP_HMAC_REG_HMAC512_KV_RD_KEY_CTRL                                                         (32'h10010600)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL                                                             (32'h600)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL_READ_EN_LOW                                                 (0)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL_READ_EN_MASK                                                (32'h1)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL_READ_ENTRY_LOW                                              (1)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL_READ_ENTRY_MASK                                             (32'h3e)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL_PCR_HASH_EXTEND_LOW                                         (6)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL_PCR_HASH_EXTEND_MASK                                        (32'h40)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL_RSVD_LOW                                                    (7)
`define HMAC_REG_HMAC512_KV_RD_KEY_CTRL_RSVD_MASK                                                   (32'hffffff80)
`define CLP_HMAC_REG_HMAC512_KV_RD_KEY_STATUS                                                       (32'h10010604)
`define HMAC_REG_HMAC512_KV_RD_KEY_STATUS                                                           (32'h604)
`define HMAC_REG_HMAC512_KV_RD_KEY_STATUS_READY_LOW                                                 (0)
`define HMAC_REG_HMAC512_KV_RD_KEY_STATUS_READY_MASK                                                (32'h1)
`define HMAC_REG_HMAC512_KV_RD_KEY_STATUS_VALID_LOW                                                 (1)
`define HMAC_REG_HMAC512_KV_RD_KEY_STATUS_VALID_MASK                                                (32'h2)
`define HMAC_REG_HMAC512_KV_RD_KEY_STATUS_ERROR_LOW                                                 (2)
`define HMAC_REG_HMAC512_KV_RD_KEY_STATUS_ERROR_MASK                                                (32'h3fc)
`define CLP_HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL                                                       (32'h10010608)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL                                                           (32'h608)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL_READ_EN_LOW                                               (0)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL_READ_EN_MASK                                              (32'h1)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL_READ_ENTRY_LOW                                            (1)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL_READ_ENTRY_MASK                                           (32'h3e)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL_PCR_HASH_EXTEND_LOW                                       (6)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL_PCR_HASH_EXTEND_MASK                                      (32'h40)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL_RSVD_LOW                                                  (7)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL_RSVD_MASK                                                 (32'hffffff80)
`define CLP_HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS                                                     (32'h1001060c)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS                                                         (32'h60c)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS_READY_LOW                                               (0)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS_READY_MASK                                              (32'h1)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS_VALID_LOW                                               (1)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS_VALID_MASK                                              (32'h2)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS_ERROR_LOW                                               (2)
`define HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS_ERROR_MASK                                              (32'h3fc)
`define CLP_HMAC_REG_HMAC512_KV_WR_CTRL                                                             (32'h10010610)
`define HMAC_REG_HMAC512_KV_WR_CTRL                                                                 (32'h610)
`define HMAC_REG_HMAC512_KV_WR_CTRL_WRITE_EN_LOW                                                    (0)
`define HMAC_REG_HMAC512_KV_WR_CTRL_WRITE_EN_MASK                                                   (32'h1)
`define HMAC_REG_HMAC512_KV_WR_CTRL_WRITE_ENTRY_LOW                                                 (1)
`define HMAC_REG_HMAC512_KV_WR_CTRL_WRITE_ENTRY_MASK                                                (32'h3e)
`define HMAC_REG_HMAC512_KV_WR_CTRL_HMAC_KEY_DEST_VALID_LOW                                         (6)
`define HMAC_REG_HMAC512_KV_WR_CTRL_HMAC_KEY_DEST_VALID_MASK                                        (32'h40)
`define HMAC_REG_HMAC512_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                       (7)
`define HMAC_REG_HMAC512_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                      (32'h80)
`define HMAC_REG_HMAC512_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_LOW                                        (8)
`define HMAC_REG_HMAC512_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_MASK                                       (32'h100)
`define HMAC_REG_HMAC512_KV_WR_CTRL_ECC_PKEY_DEST_VALID_LOW                                         (9)
`define HMAC_REG_HMAC512_KV_WR_CTRL_ECC_PKEY_DEST_VALID_MASK                                        (32'h200)
`define HMAC_REG_HMAC512_KV_WR_CTRL_ECC_SEED_DEST_VALID_LOW                                         (10)
`define HMAC_REG_HMAC512_KV_WR_CTRL_ECC_SEED_DEST_VALID_MASK                                        (32'h400)
`define HMAC_REG_HMAC512_KV_WR_CTRL_RSVD_LOW                                                        (11)
`define HMAC_REG_HMAC512_KV_WR_CTRL_RSVD_MASK                                                       (32'hfffff800)
`define CLP_HMAC_REG_HMAC512_KV_WR_STATUS                                                           (32'h10010614)
`define HMAC_REG_HMAC512_KV_WR_STATUS                                                               (32'h614)
`define HMAC_REG_HMAC512_KV_WR_STATUS_READY_LOW                                                     (0)
`define HMAC_REG_HMAC512_KV_WR_STATUS_READY_MASK                                                    (32'h1)
`define HMAC_REG_HMAC512_KV_WR_STATUS_VALID_LOW                                                     (1)
`define HMAC_REG_HMAC512_KV_WR_STATUS_VALID_MASK                                                    (32'h2)
`define HMAC_REG_HMAC512_KV_WR_STATUS_ERROR_LOW                                                     (2)
`define HMAC_REG_HMAC512_KV_WR_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_HMAC_REG_INTR_BLOCK_RF_START                                                            (32'h10010800)
`define CLP_HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                 (32'h10010800)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                     (32'h800)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                        (0)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                       (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                        (1)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                       (32'h2)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                  (32'h10010804)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                      (32'h804)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                        (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                       (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                        (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                       (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                        (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                       (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                        (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                       (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                  (32'h10010808)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                      (32'h808)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                               (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                              (32'h1001080c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                  (32'h80c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                      (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                     (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                              (32'h10010810)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                  (32'h810)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                      (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                     (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                            (32'h10010814)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                (32'h814)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                                 (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                                (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                                 (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                                (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                                 (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                                (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                                 (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                                (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                            (32'h10010818)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                (32'h818)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                         (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                        (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                (32'h1001081c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                    (32'h81c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                    (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                   (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                    (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                   (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                    (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                   (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                    (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                   (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                (32'h10010820)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                    (32'h820)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                            (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                           (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                              (32'h10010900)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                  (32'h900)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                              (32'h10010904)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                  (32'h904)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                              (32'h10010908)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                  (32'h908)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                              (32'h1001090c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                  (32'h90c)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                      (32'h10010980)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                          (32'h980)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                         (32'h10010a00)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                             (32'ha00)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                         (32'h10010a04)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                             (32'ha04)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                         (32'h10010a08)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                             (32'ha08)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                         (32'h10010a0c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                             (32'ha0c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                 (32'h10010a10)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                     (32'ha10)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                           (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                          (32'h1)
`define CLP_KV_REG_BASE_ADDR                                                                        (32'h10018000)
`define CLP_KV_REG_KEY_CTRL_0                                                                       (32'h10018000)
`define KV_REG_KEY_CTRL_0                                                                           (32'h0)
`define KV_REG_KEY_CTRL_0_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_0_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_0_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_0_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_0_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_0_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_0_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_0_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_0_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_0_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_0_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_0_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_0_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_0_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_1                                                                       (32'h10018004)
`define KV_REG_KEY_CTRL_1                                                                           (32'h4)
`define KV_REG_KEY_CTRL_1_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_1_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_1_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_1_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_1_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_1_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_1_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_1_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_1_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_1_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_1_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_1_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_1_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_1_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_2                                                                       (32'h10018008)
`define KV_REG_KEY_CTRL_2                                                                           (32'h8)
`define KV_REG_KEY_CTRL_2_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_2_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_2_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_2_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_2_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_2_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_2_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_2_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_2_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_2_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_2_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_2_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_2_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_2_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_3                                                                       (32'h1001800c)
`define KV_REG_KEY_CTRL_3                                                                           (32'hc)
`define KV_REG_KEY_CTRL_3_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_3_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_3_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_3_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_3_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_3_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_3_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_3_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_3_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_3_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_3_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_3_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_3_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_3_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_4                                                                       (32'h10018010)
`define KV_REG_KEY_CTRL_4                                                                           (32'h10)
`define KV_REG_KEY_CTRL_4_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_4_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_4_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_4_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_4_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_4_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_4_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_4_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_4_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_4_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_4_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_4_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_4_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_4_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_5                                                                       (32'h10018014)
`define KV_REG_KEY_CTRL_5                                                                           (32'h14)
`define KV_REG_KEY_CTRL_5_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_5_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_5_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_5_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_5_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_5_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_5_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_5_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_5_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_5_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_5_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_5_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_5_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_5_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_6                                                                       (32'h10018018)
`define KV_REG_KEY_CTRL_6                                                                           (32'h18)
`define KV_REG_KEY_CTRL_6_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_6_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_6_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_6_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_6_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_6_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_6_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_6_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_6_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_6_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_6_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_6_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_6_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_6_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_7                                                                       (32'h1001801c)
`define KV_REG_KEY_CTRL_7                                                                           (32'h1c)
`define KV_REG_KEY_CTRL_7_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_7_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_7_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_7_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_7_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_7_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_7_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_7_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_7_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_7_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_7_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_7_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_7_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_7_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_8                                                                       (32'h10018020)
`define KV_REG_KEY_CTRL_8                                                                           (32'h20)
`define KV_REG_KEY_CTRL_8_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_8_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_8_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_8_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_8_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_8_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_8_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_8_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_8_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_8_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_8_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_8_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_8_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_8_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_9                                                                       (32'h10018024)
`define KV_REG_KEY_CTRL_9                                                                           (32'h24)
`define KV_REG_KEY_CTRL_9_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_9_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_9_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_9_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_9_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_9_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_9_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_9_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_9_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_9_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_9_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_9_DEST_VALID_MASK                                                           (32'h1fe00)
`define KV_REG_KEY_CTRL_9_LAST_DWORD_LOW                                                            (17)
`define KV_REG_KEY_CTRL_9_LAST_DWORD_MASK                                                           (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_10                                                                      (32'h10018028)
`define KV_REG_KEY_CTRL_10                                                                          (32'h28)
`define KV_REG_KEY_CTRL_10_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_10_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_10_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_10_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_10_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_10_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_10_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_10_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_10_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_10_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_10_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_10_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_10_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_10_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_11                                                                      (32'h1001802c)
`define KV_REG_KEY_CTRL_11                                                                          (32'h2c)
`define KV_REG_KEY_CTRL_11_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_11_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_11_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_11_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_11_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_11_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_11_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_11_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_11_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_11_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_11_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_11_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_11_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_11_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_12                                                                      (32'h10018030)
`define KV_REG_KEY_CTRL_12                                                                          (32'h30)
`define KV_REG_KEY_CTRL_12_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_12_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_12_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_12_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_12_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_12_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_12_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_12_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_12_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_12_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_12_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_12_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_12_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_12_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_13                                                                      (32'h10018034)
`define KV_REG_KEY_CTRL_13                                                                          (32'h34)
`define KV_REG_KEY_CTRL_13_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_13_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_13_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_13_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_13_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_13_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_13_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_13_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_13_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_13_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_13_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_13_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_13_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_13_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_14                                                                      (32'h10018038)
`define KV_REG_KEY_CTRL_14                                                                          (32'h38)
`define KV_REG_KEY_CTRL_14_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_14_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_14_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_14_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_14_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_14_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_14_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_14_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_14_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_14_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_14_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_14_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_14_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_14_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_15                                                                      (32'h1001803c)
`define KV_REG_KEY_CTRL_15                                                                          (32'h3c)
`define KV_REG_KEY_CTRL_15_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_15_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_15_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_15_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_15_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_15_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_15_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_15_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_15_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_15_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_15_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_15_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_15_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_15_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_16                                                                      (32'h10018040)
`define KV_REG_KEY_CTRL_16                                                                          (32'h40)
`define KV_REG_KEY_CTRL_16_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_16_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_16_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_16_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_16_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_16_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_16_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_16_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_16_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_16_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_16_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_16_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_16_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_16_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_17                                                                      (32'h10018044)
`define KV_REG_KEY_CTRL_17                                                                          (32'h44)
`define KV_REG_KEY_CTRL_17_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_17_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_17_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_17_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_17_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_17_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_17_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_17_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_17_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_17_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_17_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_17_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_17_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_17_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_18                                                                      (32'h10018048)
`define KV_REG_KEY_CTRL_18                                                                          (32'h48)
`define KV_REG_KEY_CTRL_18_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_18_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_18_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_18_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_18_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_18_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_18_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_18_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_18_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_18_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_18_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_18_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_18_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_18_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_19                                                                      (32'h1001804c)
`define KV_REG_KEY_CTRL_19                                                                          (32'h4c)
`define KV_REG_KEY_CTRL_19_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_19_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_19_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_19_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_19_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_19_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_19_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_19_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_19_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_19_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_19_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_19_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_19_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_19_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_20                                                                      (32'h10018050)
`define KV_REG_KEY_CTRL_20                                                                          (32'h50)
`define KV_REG_KEY_CTRL_20_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_20_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_20_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_20_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_20_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_20_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_20_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_20_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_20_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_20_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_20_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_20_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_20_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_20_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_21                                                                      (32'h10018054)
`define KV_REG_KEY_CTRL_21                                                                          (32'h54)
`define KV_REG_KEY_CTRL_21_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_21_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_21_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_21_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_21_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_21_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_21_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_21_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_21_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_21_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_21_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_21_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_21_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_21_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_22                                                                      (32'h10018058)
`define KV_REG_KEY_CTRL_22                                                                          (32'h58)
`define KV_REG_KEY_CTRL_22_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_22_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_22_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_22_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_22_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_22_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_22_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_22_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_22_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_22_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_22_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_22_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_22_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_22_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_23                                                                      (32'h1001805c)
`define KV_REG_KEY_CTRL_23                                                                          (32'h5c)
`define KV_REG_KEY_CTRL_23_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_23_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_23_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_23_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_23_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_23_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_23_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_23_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_23_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_23_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_23_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_23_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_23_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_23_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_24                                                                      (32'h10018060)
`define KV_REG_KEY_CTRL_24                                                                          (32'h60)
`define KV_REG_KEY_CTRL_24_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_24_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_24_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_24_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_24_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_24_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_24_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_24_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_24_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_24_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_24_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_24_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_24_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_24_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_25                                                                      (32'h10018064)
`define KV_REG_KEY_CTRL_25                                                                          (32'h64)
`define KV_REG_KEY_CTRL_25_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_25_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_25_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_25_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_25_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_25_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_25_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_25_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_25_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_25_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_25_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_25_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_25_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_25_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_26                                                                      (32'h10018068)
`define KV_REG_KEY_CTRL_26                                                                          (32'h68)
`define KV_REG_KEY_CTRL_26_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_26_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_26_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_26_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_26_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_26_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_26_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_26_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_26_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_26_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_26_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_26_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_26_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_26_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_27                                                                      (32'h1001806c)
`define KV_REG_KEY_CTRL_27                                                                          (32'h6c)
`define KV_REG_KEY_CTRL_27_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_27_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_27_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_27_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_27_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_27_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_27_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_27_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_27_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_27_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_27_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_27_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_27_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_27_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_28                                                                      (32'h10018070)
`define KV_REG_KEY_CTRL_28                                                                          (32'h70)
`define KV_REG_KEY_CTRL_28_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_28_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_28_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_28_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_28_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_28_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_28_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_28_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_28_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_28_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_28_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_28_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_28_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_28_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_29                                                                      (32'h10018074)
`define KV_REG_KEY_CTRL_29                                                                          (32'h74)
`define KV_REG_KEY_CTRL_29_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_29_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_29_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_29_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_29_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_29_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_29_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_29_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_29_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_29_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_29_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_29_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_29_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_29_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_30                                                                      (32'h10018078)
`define KV_REG_KEY_CTRL_30                                                                          (32'h78)
`define KV_REG_KEY_CTRL_30_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_30_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_30_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_30_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_30_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_30_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_30_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_30_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_30_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_30_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_30_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_30_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_30_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_30_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_CTRL_31                                                                      (32'h1001807c)
`define KV_REG_KEY_CTRL_31                                                                          (32'h7c)
`define KV_REG_KEY_CTRL_31_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_31_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_31_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_31_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_31_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_31_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_31_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_31_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_31_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_31_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_31_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_31_DEST_VALID_MASK                                                          (32'h1fe00)
`define KV_REG_KEY_CTRL_31_LAST_DWORD_LOW                                                           (17)
`define KV_REG_KEY_CTRL_31_LAST_DWORD_MASK                                                          (32'h1e0000)
`define CLP_KV_REG_KEY_ENTRY_0_0                                                                    (32'h10018600)
`define KV_REG_KEY_ENTRY_0_0                                                                        (32'h600)
`define CLP_KV_REG_KEY_ENTRY_0_1                                                                    (32'h10018604)
`define KV_REG_KEY_ENTRY_0_1                                                                        (32'h604)
`define CLP_KV_REG_KEY_ENTRY_0_2                                                                    (32'h10018608)
`define KV_REG_KEY_ENTRY_0_2                                                                        (32'h608)
`define CLP_KV_REG_KEY_ENTRY_0_3                                                                    (32'h1001860c)
`define KV_REG_KEY_ENTRY_0_3                                                                        (32'h60c)
`define CLP_KV_REG_KEY_ENTRY_0_4                                                                    (32'h10018610)
`define KV_REG_KEY_ENTRY_0_4                                                                        (32'h610)
`define CLP_KV_REG_KEY_ENTRY_0_5                                                                    (32'h10018614)
`define KV_REG_KEY_ENTRY_0_5                                                                        (32'h614)
`define CLP_KV_REG_KEY_ENTRY_0_6                                                                    (32'h10018618)
`define KV_REG_KEY_ENTRY_0_6                                                                        (32'h618)
`define CLP_KV_REG_KEY_ENTRY_0_7                                                                    (32'h1001861c)
`define KV_REG_KEY_ENTRY_0_7                                                                        (32'h61c)
`define CLP_KV_REG_KEY_ENTRY_0_8                                                                    (32'h10018620)
`define KV_REG_KEY_ENTRY_0_8                                                                        (32'h620)
`define CLP_KV_REG_KEY_ENTRY_0_9                                                                    (32'h10018624)
`define KV_REG_KEY_ENTRY_0_9                                                                        (32'h624)
`define CLP_KV_REG_KEY_ENTRY_0_10                                                                   (32'h10018628)
`define KV_REG_KEY_ENTRY_0_10                                                                       (32'h628)
`define CLP_KV_REG_KEY_ENTRY_0_11                                                                   (32'h1001862c)
`define KV_REG_KEY_ENTRY_0_11                                                                       (32'h62c)
`define CLP_KV_REG_KEY_ENTRY_1_0                                                                    (32'h10018630)
`define KV_REG_KEY_ENTRY_1_0                                                                        (32'h630)
`define CLP_KV_REG_KEY_ENTRY_1_1                                                                    (32'h10018634)
`define KV_REG_KEY_ENTRY_1_1                                                                        (32'h634)
`define CLP_KV_REG_KEY_ENTRY_1_2                                                                    (32'h10018638)
`define KV_REG_KEY_ENTRY_1_2                                                                        (32'h638)
`define CLP_KV_REG_KEY_ENTRY_1_3                                                                    (32'h1001863c)
`define KV_REG_KEY_ENTRY_1_3                                                                        (32'h63c)
`define CLP_KV_REG_KEY_ENTRY_1_4                                                                    (32'h10018640)
`define KV_REG_KEY_ENTRY_1_4                                                                        (32'h640)
`define CLP_KV_REG_KEY_ENTRY_1_5                                                                    (32'h10018644)
`define KV_REG_KEY_ENTRY_1_5                                                                        (32'h644)
`define CLP_KV_REG_KEY_ENTRY_1_6                                                                    (32'h10018648)
`define KV_REG_KEY_ENTRY_1_6                                                                        (32'h648)
`define CLP_KV_REG_KEY_ENTRY_1_7                                                                    (32'h1001864c)
`define KV_REG_KEY_ENTRY_1_7                                                                        (32'h64c)
`define CLP_KV_REG_KEY_ENTRY_1_8                                                                    (32'h10018650)
`define KV_REG_KEY_ENTRY_1_8                                                                        (32'h650)
`define CLP_KV_REG_KEY_ENTRY_1_9                                                                    (32'h10018654)
`define KV_REG_KEY_ENTRY_1_9                                                                        (32'h654)
`define CLP_KV_REG_KEY_ENTRY_1_10                                                                   (32'h10018658)
`define KV_REG_KEY_ENTRY_1_10                                                                       (32'h658)
`define CLP_KV_REG_KEY_ENTRY_1_11                                                                   (32'h1001865c)
`define KV_REG_KEY_ENTRY_1_11                                                                       (32'h65c)
`define CLP_KV_REG_KEY_ENTRY_2_0                                                                    (32'h10018660)
`define KV_REG_KEY_ENTRY_2_0                                                                        (32'h660)
`define CLP_KV_REG_KEY_ENTRY_2_1                                                                    (32'h10018664)
`define KV_REG_KEY_ENTRY_2_1                                                                        (32'h664)
`define CLP_KV_REG_KEY_ENTRY_2_2                                                                    (32'h10018668)
`define KV_REG_KEY_ENTRY_2_2                                                                        (32'h668)
`define CLP_KV_REG_KEY_ENTRY_2_3                                                                    (32'h1001866c)
`define KV_REG_KEY_ENTRY_2_3                                                                        (32'h66c)
`define CLP_KV_REG_KEY_ENTRY_2_4                                                                    (32'h10018670)
`define KV_REG_KEY_ENTRY_2_4                                                                        (32'h670)
`define CLP_KV_REG_KEY_ENTRY_2_5                                                                    (32'h10018674)
`define KV_REG_KEY_ENTRY_2_5                                                                        (32'h674)
`define CLP_KV_REG_KEY_ENTRY_2_6                                                                    (32'h10018678)
`define KV_REG_KEY_ENTRY_2_6                                                                        (32'h678)
`define CLP_KV_REG_KEY_ENTRY_2_7                                                                    (32'h1001867c)
`define KV_REG_KEY_ENTRY_2_7                                                                        (32'h67c)
`define CLP_KV_REG_KEY_ENTRY_2_8                                                                    (32'h10018680)
`define KV_REG_KEY_ENTRY_2_8                                                                        (32'h680)
`define CLP_KV_REG_KEY_ENTRY_2_9                                                                    (32'h10018684)
`define KV_REG_KEY_ENTRY_2_9                                                                        (32'h684)
`define CLP_KV_REG_KEY_ENTRY_2_10                                                                   (32'h10018688)
`define KV_REG_KEY_ENTRY_2_10                                                                       (32'h688)
`define CLP_KV_REG_KEY_ENTRY_2_11                                                                   (32'h1001868c)
`define KV_REG_KEY_ENTRY_2_11                                                                       (32'h68c)
`define CLP_KV_REG_KEY_ENTRY_3_0                                                                    (32'h10018690)
`define KV_REG_KEY_ENTRY_3_0                                                                        (32'h690)
`define CLP_KV_REG_KEY_ENTRY_3_1                                                                    (32'h10018694)
`define KV_REG_KEY_ENTRY_3_1                                                                        (32'h694)
`define CLP_KV_REG_KEY_ENTRY_3_2                                                                    (32'h10018698)
`define KV_REG_KEY_ENTRY_3_2                                                                        (32'h698)
`define CLP_KV_REG_KEY_ENTRY_3_3                                                                    (32'h1001869c)
`define KV_REG_KEY_ENTRY_3_3                                                                        (32'h69c)
`define CLP_KV_REG_KEY_ENTRY_3_4                                                                    (32'h100186a0)
`define KV_REG_KEY_ENTRY_3_4                                                                        (32'h6a0)
`define CLP_KV_REG_KEY_ENTRY_3_5                                                                    (32'h100186a4)
`define KV_REG_KEY_ENTRY_3_5                                                                        (32'h6a4)
`define CLP_KV_REG_KEY_ENTRY_3_6                                                                    (32'h100186a8)
`define KV_REG_KEY_ENTRY_3_6                                                                        (32'h6a8)
`define CLP_KV_REG_KEY_ENTRY_3_7                                                                    (32'h100186ac)
`define KV_REG_KEY_ENTRY_3_7                                                                        (32'h6ac)
`define CLP_KV_REG_KEY_ENTRY_3_8                                                                    (32'h100186b0)
`define KV_REG_KEY_ENTRY_3_8                                                                        (32'h6b0)
`define CLP_KV_REG_KEY_ENTRY_3_9                                                                    (32'h100186b4)
`define KV_REG_KEY_ENTRY_3_9                                                                        (32'h6b4)
`define CLP_KV_REG_KEY_ENTRY_3_10                                                                   (32'h100186b8)
`define KV_REG_KEY_ENTRY_3_10                                                                       (32'h6b8)
`define CLP_KV_REG_KEY_ENTRY_3_11                                                                   (32'h100186bc)
`define KV_REG_KEY_ENTRY_3_11                                                                       (32'h6bc)
`define CLP_KV_REG_KEY_ENTRY_4_0                                                                    (32'h100186c0)
`define KV_REG_KEY_ENTRY_4_0                                                                        (32'h6c0)
`define CLP_KV_REG_KEY_ENTRY_4_1                                                                    (32'h100186c4)
`define KV_REG_KEY_ENTRY_4_1                                                                        (32'h6c4)
`define CLP_KV_REG_KEY_ENTRY_4_2                                                                    (32'h100186c8)
`define KV_REG_KEY_ENTRY_4_2                                                                        (32'h6c8)
`define CLP_KV_REG_KEY_ENTRY_4_3                                                                    (32'h100186cc)
`define KV_REG_KEY_ENTRY_4_3                                                                        (32'h6cc)
`define CLP_KV_REG_KEY_ENTRY_4_4                                                                    (32'h100186d0)
`define KV_REG_KEY_ENTRY_4_4                                                                        (32'h6d0)
`define CLP_KV_REG_KEY_ENTRY_4_5                                                                    (32'h100186d4)
`define KV_REG_KEY_ENTRY_4_5                                                                        (32'h6d4)
`define CLP_KV_REG_KEY_ENTRY_4_6                                                                    (32'h100186d8)
`define KV_REG_KEY_ENTRY_4_6                                                                        (32'h6d8)
`define CLP_KV_REG_KEY_ENTRY_4_7                                                                    (32'h100186dc)
`define KV_REG_KEY_ENTRY_4_7                                                                        (32'h6dc)
`define CLP_KV_REG_KEY_ENTRY_4_8                                                                    (32'h100186e0)
`define KV_REG_KEY_ENTRY_4_8                                                                        (32'h6e0)
`define CLP_KV_REG_KEY_ENTRY_4_9                                                                    (32'h100186e4)
`define KV_REG_KEY_ENTRY_4_9                                                                        (32'h6e4)
`define CLP_KV_REG_KEY_ENTRY_4_10                                                                   (32'h100186e8)
`define KV_REG_KEY_ENTRY_4_10                                                                       (32'h6e8)
`define CLP_KV_REG_KEY_ENTRY_4_11                                                                   (32'h100186ec)
`define KV_REG_KEY_ENTRY_4_11                                                                       (32'h6ec)
`define CLP_KV_REG_KEY_ENTRY_5_0                                                                    (32'h100186f0)
`define KV_REG_KEY_ENTRY_5_0                                                                        (32'h6f0)
`define CLP_KV_REG_KEY_ENTRY_5_1                                                                    (32'h100186f4)
`define KV_REG_KEY_ENTRY_5_1                                                                        (32'h6f4)
`define CLP_KV_REG_KEY_ENTRY_5_2                                                                    (32'h100186f8)
`define KV_REG_KEY_ENTRY_5_2                                                                        (32'h6f8)
`define CLP_KV_REG_KEY_ENTRY_5_3                                                                    (32'h100186fc)
`define KV_REG_KEY_ENTRY_5_3                                                                        (32'h6fc)
`define CLP_KV_REG_KEY_ENTRY_5_4                                                                    (32'h10018700)
`define KV_REG_KEY_ENTRY_5_4                                                                        (32'h700)
`define CLP_KV_REG_KEY_ENTRY_5_5                                                                    (32'h10018704)
`define KV_REG_KEY_ENTRY_5_5                                                                        (32'h704)
`define CLP_KV_REG_KEY_ENTRY_5_6                                                                    (32'h10018708)
`define KV_REG_KEY_ENTRY_5_6                                                                        (32'h708)
`define CLP_KV_REG_KEY_ENTRY_5_7                                                                    (32'h1001870c)
`define KV_REG_KEY_ENTRY_5_7                                                                        (32'h70c)
`define CLP_KV_REG_KEY_ENTRY_5_8                                                                    (32'h10018710)
`define KV_REG_KEY_ENTRY_5_8                                                                        (32'h710)
`define CLP_KV_REG_KEY_ENTRY_5_9                                                                    (32'h10018714)
`define KV_REG_KEY_ENTRY_5_9                                                                        (32'h714)
`define CLP_KV_REG_KEY_ENTRY_5_10                                                                   (32'h10018718)
`define KV_REG_KEY_ENTRY_5_10                                                                       (32'h718)
`define CLP_KV_REG_KEY_ENTRY_5_11                                                                   (32'h1001871c)
`define KV_REG_KEY_ENTRY_5_11                                                                       (32'h71c)
`define CLP_KV_REG_KEY_ENTRY_6_0                                                                    (32'h10018720)
`define KV_REG_KEY_ENTRY_6_0                                                                        (32'h720)
`define CLP_KV_REG_KEY_ENTRY_6_1                                                                    (32'h10018724)
`define KV_REG_KEY_ENTRY_6_1                                                                        (32'h724)
`define CLP_KV_REG_KEY_ENTRY_6_2                                                                    (32'h10018728)
`define KV_REG_KEY_ENTRY_6_2                                                                        (32'h728)
`define CLP_KV_REG_KEY_ENTRY_6_3                                                                    (32'h1001872c)
`define KV_REG_KEY_ENTRY_6_3                                                                        (32'h72c)
`define CLP_KV_REG_KEY_ENTRY_6_4                                                                    (32'h10018730)
`define KV_REG_KEY_ENTRY_6_4                                                                        (32'h730)
`define CLP_KV_REG_KEY_ENTRY_6_5                                                                    (32'h10018734)
`define KV_REG_KEY_ENTRY_6_5                                                                        (32'h734)
`define CLP_KV_REG_KEY_ENTRY_6_6                                                                    (32'h10018738)
`define KV_REG_KEY_ENTRY_6_6                                                                        (32'h738)
`define CLP_KV_REG_KEY_ENTRY_6_7                                                                    (32'h1001873c)
`define KV_REG_KEY_ENTRY_6_7                                                                        (32'h73c)
`define CLP_KV_REG_KEY_ENTRY_6_8                                                                    (32'h10018740)
`define KV_REG_KEY_ENTRY_6_8                                                                        (32'h740)
`define CLP_KV_REG_KEY_ENTRY_6_9                                                                    (32'h10018744)
`define KV_REG_KEY_ENTRY_6_9                                                                        (32'h744)
`define CLP_KV_REG_KEY_ENTRY_6_10                                                                   (32'h10018748)
`define KV_REG_KEY_ENTRY_6_10                                                                       (32'h748)
`define CLP_KV_REG_KEY_ENTRY_6_11                                                                   (32'h1001874c)
`define KV_REG_KEY_ENTRY_6_11                                                                       (32'h74c)
`define CLP_KV_REG_KEY_ENTRY_7_0                                                                    (32'h10018750)
`define KV_REG_KEY_ENTRY_7_0                                                                        (32'h750)
`define CLP_KV_REG_KEY_ENTRY_7_1                                                                    (32'h10018754)
`define KV_REG_KEY_ENTRY_7_1                                                                        (32'h754)
`define CLP_KV_REG_KEY_ENTRY_7_2                                                                    (32'h10018758)
`define KV_REG_KEY_ENTRY_7_2                                                                        (32'h758)
`define CLP_KV_REG_KEY_ENTRY_7_3                                                                    (32'h1001875c)
`define KV_REG_KEY_ENTRY_7_3                                                                        (32'h75c)
`define CLP_KV_REG_KEY_ENTRY_7_4                                                                    (32'h10018760)
`define KV_REG_KEY_ENTRY_7_4                                                                        (32'h760)
`define CLP_KV_REG_KEY_ENTRY_7_5                                                                    (32'h10018764)
`define KV_REG_KEY_ENTRY_7_5                                                                        (32'h764)
`define CLP_KV_REG_KEY_ENTRY_7_6                                                                    (32'h10018768)
`define KV_REG_KEY_ENTRY_7_6                                                                        (32'h768)
`define CLP_KV_REG_KEY_ENTRY_7_7                                                                    (32'h1001876c)
`define KV_REG_KEY_ENTRY_7_7                                                                        (32'h76c)
`define CLP_KV_REG_KEY_ENTRY_7_8                                                                    (32'h10018770)
`define KV_REG_KEY_ENTRY_7_8                                                                        (32'h770)
`define CLP_KV_REG_KEY_ENTRY_7_9                                                                    (32'h10018774)
`define KV_REG_KEY_ENTRY_7_9                                                                        (32'h774)
`define CLP_KV_REG_KEY_ENTRY_7_10                                                                   (32'h10018778)
`define KV_REG_KEY_ENTRY_7_10                                                                       (32'h778)
`define CLP_KV_REG_KEY_ENTRY_7_11                                                                   (32'h1001877c)
`define KV_REG_KEY_ENTRY_7_11                                                                       (32'h77c)
`define CLP_KV_REG_KEY_ENTRY_8_0                                                                    (32'h10018780)
`define KV_REG_KEY_ENTRY_8_0                                                                        (32'h780)
`define CLP_KV_REG_KEY_ENTRY_8_1                                                                    (32'h10018784)
`define KV_REG_KEY_ENTRY_8_1                                                                        (32'h784)
`define CLP_KV_REG_KEY_ENTRY_8_2                                                                    (32'h10018788)
`define KV_REG_KEY_ENTRY_8_2                                                                        (32'h788)
`define CLP_KV_REG_KEY_ENTRY_8_3                                                                    (32'h1001878c)
`define KV_REG_KEY_ENTRY_8_3                                                                        (32'h78c)
`define CLP_KV_REG_KEY_ENTRY_8_4                                                                    (32'h10018790)
`define KV_REG_KEY_ENTRY_8_4                                                                        (32'h790)
`define CLP_KV_REG_KEY_ENTRY_8_5                                                                    (32'h10018794)
`define KV_REG_KEY_ENTRY_8_5                                                                        (32'h794)
`define CLP_KV_REG_KEY_ENTRY_8_6                                                                    (32'h10018798)
`define KV_REG_KEY_ENTRY_8_6                                                                        (32'h798)
`define CLP_KV_REG_KEY_ENTRY_8_7                                                                    (32'h1001879c)
`define KV_REG_KEY_ENTRY_8_7                                                                        (32'h79c)
`define CLP_KV_REG_KEY_ENTRY_8_8                                                                    (32'h100187a0)
`define KV_REG_KEY_ENTRY_8_8                                                                        (32'h7a0)
`define CLP_KV_REG_KEY_ENTRY_8_9                                                                    (32'h100187a4)
`define KV_REG_KEY_ENTRY_8_9                                                                        (32'h7a4)
`define CLP_KV_REG_KEY_ENTRY_8_10                                                                   (32'h100187a8)
`define KV_REG_KEY_ENTRY_8_10                                                                       (32'h7a8)
`define CLP_KV_REG_KEY_ENTRY_8_11                                                                   (32'h100187ac)
`define KV_REG_KEY_ENTRY_8_11                                                                       (32'h7ac)
`define CLP_KV_REG_KEY_ENTRY_9_0                                                                    (32'h100187b0)
`define KV_REG_KEY_ENTRY_9_0                                                                        (32'h7b0)
`define CLP_KV_REG_KEY_ENTRY_9_1                                                                    (32'h100187b4)
`define KV_REG_KEY_ENTRY_9_1                                                                        (32'h7b4)
`define CLP_KV_REG_KEY_ENTRY_9_2                                                                    (32'h100187b8)
`define KV_REG_KEY_ENTRY_9_2                                                                        (32'h7b8)
`define CLP_KV_REG_KEY_ENTRY_9_3                                                                    (32'h100187bc)
`define KV_REG_KEY_ENTRY_9_3                                                                        (32'h7bc)
`define CLP_KV_REG_KEY_ENTRY_9_4                                                                    (32'h100187c0)
`define KV_REG_KEY_ENTRY_9_4                                                                        (32'h7c0)
`define CLP_KV_REG_KEY_ENTRY_9_5                                                                    (32'h100187c4)
`define KV_REG_KEY_ENTRY_9_5                                                                        (32'h7c4)
`define CLP_KV_REG_KEY_ENTRY_9_6                                                                    (32'h100187c8)
`define KV_REG_KEY_ENTRY_9_6                                                                        (32'h7c8)
`define CLP_KV_REG_KEY_ENTRY_9_7                                                                    (32'h100187cc)
`define KV_REG_KEY_ENTRY_9_7                                                                        (32'h7cc)
`define CLP_KV_REG_KEY_ENTRY_9_8                                                                    (32'h100187d0)
`define KV_REG_KEY_ENTRY_9_8                                                                        (32'h7d0)
`define CLP_KV_REG_KEY_ENTRY_9_9                                                                    (32'h100187d4)
`define KV_REG_KEY_ENTRY_9_9                                                                        (32'h7d4)
`define CLP_KV_REG_KEY_ENTRY_9_10                                                                   (32'h100187d8)
`define KV_REG_KEY_ENTRY_9_10                                                                       (32'h7d8)
`define CLP_KV_REG_KEY_ENTRY_9_11                                                                   (32'h100187dc)
`define KV_REG_KEY_ENTRY_9_11                                                                       (32'h7dc)
`define CLP_KV_REG_KEY_ENTRY_10_0                                                                   (32'h100187e0)
`define KV_REG_KEY_ENTRY_10_0                                                                       (32'h7e0)
`define CLP_KV_REG_KEY_ENTRY_10_1                                                                   (32'h100187e4)
`define KV_REG_KEY_ENTRY_10_1                                                                       (32'h7e4)
`define CLP_KV_REG_KEY_ENTRY_10_2                                                                   (32'h100187e8)
`define KV_REG_KEY_ENTRY_10_2                                                                       (32'h7e8)
`define CLP_KV_REG_KEY_ENTRY_10_3                                                                   (32'h100187ec)
`define KV_REG_KEY_ENTRY_10_3                                                                       (32'h7ec)
`define CLP_KV_REG_KEY_ENTRY_10_4                                                                   (32'h100187f0)
`define KV_REG_KEY_ENTRY_10_4                                                                       (32'h7f0)
`define CLP_KV_REG_KEY_ENTRY_10_5                                                                   (32'h100187f4)
`define KV_REG_KEY_ENTRY_10_5                                                                       (32'h7f4)
`define CLP_KV_REG_KEY_ENTRY_10_6                                                                   (32'h100187f8)
`define KV_REG_KEY_ENTRY_10_6                                                                       (32'h7f8)
`define CLP_KV_REG_KEY_ENTRY_10_7                                                                   (32'h100187fc)
`define KV_REG_KEY_ENTRY_10_7                                                                       (32'h7fc)
`define CLP_KV_REG_KEY_ENTRY_10_8                                                                   (32'h10018800)
`define KV_REG_KEY_ENTRY_10_8                                                                       (32'h800)
`define CLP_KV_REG_KEY_ENTRY_10_9                                                                   (32'h10018804)
`define KV_REG_KEY_ENTRY_10_9                                                                       (32'h804)
`define CLP_KV_REG_KEY_ENTRY_10_10                                                                  (32'h10018808)
`define KV_REG_KEY_ENTRY_10_10                                                                      (32'h808)
`define CLP_KV_REG_KEY_ENTRY_10_11                                                                  (32'h1001880c)
`define KV_REG_KEY_ENTRY_10_11                                                                      (32'h80c)
`define CLP_KV_REG_KEY_ENTRY_11_0                                                                   (32'h10018810)
`define KV_REG_KEY_ENTRY_11_0                                                                       (32'h810)
`define CLP_KV_REG_KEY_ENTRY_11_1                                                                   (32'h10018814)
`define KV_REG_KEY_ENTRY_11_1                                                                       (32'h814)
`define CLP_KV_REG_KEY_ENTRY_11_2                                                                   (32'h10018818)
`define KV_REG_KEY_ENTRY_11_2                                                                       (32'h818)
`define CLP_KV_REG_KEY_ENTRY_11_3                                                                   (32'h1001881c)
`define KV_REG_KEY_ENTRY_11_3                                                                       (32'h81c)
`define CLP_KV_REG_KEY_ENTRY_11_4                                                                   (32'h10018820)
`define KV_REG_KEY_ENTRY_11_4                                                                       (32'h820)
`define CLP_KV_REG_KEY_ENTRY_11_5                                                                   (32'h10018824)
`define KV_REG_KEY_ENTRY_11_5                                                                       (32'h824)
`define CLP_KV_REG_KEY_ENTRY_11_6                                                                   (32'h10018828)
`define KV_REG_KEY_ENTRY_11_6                                                                       (32'h828)
`define CLP_KV_REG_KEY_ENTRY_11_7                                                                   (32'h1001882c)
`define KV_REG_KEY_ENTRY_11_7                                                                       (32'h82c)
`define CLP_KV_REG_KEY_ENTRY_11_8                                                                   (32'h10018830)
`define KV_REG_KEY_ENTRY_11_8                                                                       (32'h830)
`define CLP_KV_REG_KEY_ENTRY_11_9                                                                   (32'h10018834)
`define KV_REG_KEY_ENTRY_11_9                                                                       (32'h834)
`define CLP_KV_REG_KEY_ENTRY_11_10                                                                  (32'h10018838)
`define KV_REG_KEY_ENTRY_11_10                                                                      (32'h838)
`define CLP_KV_REG_KEY_ENTRY_11_11                                                                  (32'h1001883c)
`define KV_REG_KEY_ENTRY_11_11                                                                      (32'h83c)
`define CLP_KV_REG_KEY_ENTRY_12_0                                                                   (32'h10018840)
`define KV_REG_KEY_ENTRY_12_0                                                                       (32'h840)
`define CLP_KV_REG_KEY_ENTRY_12_1                                                                   (32'h10018844)
`define KV_REG_KEY_ENTRY_12_1                                                                       (32'h844)
`define CLP_KV_REG_KEY_ENTRY_12_2                                                                   (32'h10018848)
`define KV_REG_KEY_ENTRY_12_2                                                                       (32'h848)
`define CLP_KV_REG_KEY_ENTRY_12_3                                                                   (32'h1001884c)
`define KV_REG_KEY_ENTRY_12_3                                                                       (32'h84c)
`define CLP_KV_REG_KEY_ENTRY_12_4                                                                   (32'h10018850)
`define KV_REG_KEY_ENTRY_12_4                                                                       (32'h850)
`define CLP_KV_REG_KEY_ENTRY_12_5                                                                   (32'h10018854)
`define KV_REG_KEY_ENTRY_12_5                                                                       (32'h854)
`define CLP_KV_REG_KEY_ENTRY_12_6                                                                   (32'h10018858)
`define KV_REG_KEY_ENTRY_12_6                                                                       (32'h858)
`define CLP_KV_REG_KEY_ENTRY_12_7                                                                   (32'h1001885c)
`define KV_REG_KEY_ENTRY_12_7                                                                       (32'h85c)
`define CLP_KV_REG_KEY_ENTRY_12_8                                                                   (32'h10018860)
`define KV_REG_KEY_ENTRY_12_8                                                                       (32'h860)
`define CLP_KV_REG_KEY_ENTRY_12_9                                                                   (32'h10018864)
`define KV_REG_KEY_ENTRY_12_9                                                                       (32'h864)
`define CLP_KV_REG_KEY_ENTRY_12_10                                                                  (32'h10018868)
`define KV_REG_KEY_ENTRY_12_10                                                                      (32'h868)
`define CLP_KV_REG_KEY_ENTRY_12_11                                                                  (32'h1001886c)
`define KV_REG_KEY_ENTRY_12_11                                                                      (32'h86c)
`define CLP_KV_REG_KEY_ENTRY_13_0                                                                   (32'h10018870)
`define KV_REG_KEY_ENTRY_13_0                                                                       (32'h870)
`define CLP_KV_REG_KEY_ENTRY_13_1                                                                   (32'h10018874)
`define KV_REG_KEY_ENTRY_13_1                                                                       (32'h874)
`define CLP_KV_REG_KEY_ENTRY_13_2                                                                   (32'h10018878)
`define KV_REG_KEY_ENTRY_13_2                                                                       (32'h878)
`define CLP_KV_REG_KEY_ENTRY_13_3                                                                   (32'h1001887c)
`define KV_REG_KEY_ENTRY_13_3                                                                       (32'h87c)
`define CLP_KV_REG_KEY_ENTRY_13_4                                                                   (32'h10018880)
`define KV_REG_KEY_ENTRY_13_4                                                                       (32'h880)
`define CLP_KV_REG_KEY_ENTRY_13_5                                                                   (32'h10018884)
`define KV_REG_KEY_ENTRY_13_5                                                                       (32'h884)
`define CLP_KV_REG_KEY_ENTRY_13_6                                                                   (32'h10018888)
`define KV_REG_KEY_ENTRY_13_6                                                                       (32'h888)
`define CLP_KV_REG_KEY_ENTRY_13_7                                                                   (32'h1001888c)
`define KV_REG_KEY_ENTRY_13_7                                                                       (32'h88c)
`define CLP_KV_REG_KEY_ENTRY_13_8                                                                   (32'h10018890)
`define KV_REG_KEY_ENTRY_13_8                                                                       (32'h890)
`define CLP_KV_REG_KEY_ENTRY_13_9                                                                   (32'h10018894)
`define KV_REG_KEY_ENTRY_13_9                                                                       (32'h894)
`define CLP_KV_REG_KEY_ENTRY_13_10                                                                  (32'h10018898)
`define KV_REG_KEY_ENTRY_13_10                                                                      (32'h898)
`define CLP_KV_REG_KEY_ENTRY_13_11                                                                  (32'h1001889c)
`define KV_REG_KEY_ENTRY_13_11                                                                      (32'h89c)
`define CLP_KV_REG_KEY_ENTRY_14_0                                                                   (32'h100188a0)
`define KV_REG_KEY_ENTRY_14_0                                                                       (32'h8a0)
`define CLP_KV_REG_KEY_ENTRY_14_1                                                                   (32'h100188a4)
`define KV_REG_KEY_ENTRY_14_1                                                                       (32'h8a4)
`define CLP_KV_REG_KEY_ENTRY_14_2                                                                   (32'h100188a8)
`define KV_REG_KEY_ENTRY_14_2                                                                       (32'h8a8)
`define CLP_KV_REG_KEY_ENTRY_14_3                                                                   (32'h100188ac)
`define KV_REG_KEY_ENTRY_14_3                                                                       (32'h8ac)
`define CLP_KV_REG_KEY_ENTRY_14_4                                                                   (32'h100188b0)
`define KV_REG_KEY_ENTRY_14_4                                                                       (32'h8b0)
`define CLP_KV_REG_KEY_ENTRY_14_5                                                                   (32'h100188b4)
`define KV_REG_KEY_ENTRY_14_5                                                                       (32'h8b4)
`define CLP_KV_REG_KEY_ENTRY_14_6                                                                   (32'h100188b8)
`define KV_REG_KEY_ENTRY_14_6                                                                       (32'h8b8)
`define CLP_KV_REG_KEY_ENTRY_14_7                                                                   (32'h100188bc)
`define KV_REG_KEY_ENTRY_14_7                                                                       (32'h8bc)
`define CLP_KV_REG_KEY_ENTRY_14_8                                                                   (32'h100188c0)
`define KV_REG_KEY_ENTRY_14_8                                                                       (32'h8c0)
`define CLP_KV_REG_KEY_ENTRY_14_9                                                                   (32'h100188c4)
`define KV_REG_KEY_ENTRY_14_9                                                                       (32'h8c4)
`define CLP_KV_REG_KEY_ENTRY_14_10                                                                  (32'h100188c8)
`define KV_REG_KEY_ENTRY_14_10                                                                      (32'h8c8)
`define CLP_KV_REG_KEY_ENTRY_14_11                                                                  (32'h100188cc)
`define KV_REG_KEY_ENTRY_14_11                                                                      (32'h8cc)
`define CLP_KV_REG_KEY_ENTRY_15_0                                                                   (32'h100188d0)
`define KV_REG_KEY_ENTRY_15_0                                                                       (32'h8d0)
`define CLP_KV_REG_KEY_ENTRY_15_1                                                                   (32'h100188d4)
`define KV_REG_KEY_ENTRY_15_1                                                                       (32'h8d4)
`define CLP_KV_REG_KEY_ENTRY_15_2                                                                   (32'h100188d8)
`define KV_REG_KEY_ENTRY_15_2                                                                       (32'h8d8)
`define CLP_KV_REG_KEY_ENTRY_15_3                                                                   (32'h100188dc)
`define KV_REG_KEY_ENTRY_15_3                                                                       (32'h8dc)
`define CLP_KV_REG_KEY_ENTRY_15_4                                                                   (32'h100188e0)
`define KV_REG_KEY_ENTRY_15_4                                                                       (32'h8e0)
`define CLP_KV_REG_KEY_ENTRY_15_5                                                                   (32'h100188e4)
`define KV_REG_KEY_ENTRY_15_5                                                                       (32'h8e4)
`define CLP_KV_REG_KEY_ENTRY_15_6                                                                   (32'h100188e8)
`define KV_REG_KEY_ENTRY_15_6                                                                       (32'h8e8)
`define CLP_KV_REG_KEY_ENTRY_15_7                                                                   (32'h100188ec)
`define KV_REG_KEY_ENTRY_15_7                                                                       (32'h8ec)
`define CLP_KV_REG_KEY_ENTRY_15_8                                                                   (32'h100188f0)
`define KV_REG_KEY_ENTRY_15_8                                                                       (32'h8f0)
`define CLP_KV_REG_KEY_ENTRY_15_9                                                                   (32'h100188f4)
`define KV_REG_KEY_ENTRY_15_9                                                                       (32'h8f4)
`define CLP_KV_REG_KEY_ENTRY_15_10                                                                  (32'h100188f8)
`define KV_REG_KEY_ENTRY_15_10                                                                      (32'h8f8)
`define CLP_KV_REG_KEY_ENTRY_15_11                                                                  (32'h100188fc)
`define KV_REG_KEY_ENTRY_15_11                                                                      (32'h8fc)
`define CLP_KV_REG_KEY_ENTRY_16_0                                                                   (32'h10018900)
`define KV_REG_KEY_ENTRY_16_0                                                                       (32'h900)
`define CLP_KV_REG_KEY_ENTRY_16_1                                                                   (32'h10018904)
`define KV_REG_KEY_ENTRY_16_1                                                                       (32'h904)
`define CLP_KV_REG_KEY_ENTRY_16_2                                                                   (32'h10018908)
`define KV_REG_KEY_ENTRY_16_2                                                                       (32'h908)
`define CLP_KV_REG_KEY_ENTRY_16_3                                                                   (32'h1001890c)
`define KV_REG_KEY_ENTRY_16_3                                                                       (32'h90c)
`define CLP_KV_REG_KEY_ENTRY_16_4                                                                   (32'h10018910)
`define KV_REG_KEY_ENTRY_16_4                                                                       (32'h910)
`define CLP_KV_REG_KEY_ENTRY_16_5                                                                   (32'h10018914)
`define KV_REG_KEY_ENTRY_16_5                                                                       (32'h914)
`define CLP_KV_REG_KEY_ENTRY_16_6                                                                   (32'h10018918)
`define KV_REG_KEY_ENTRY_16_6                                                                       (32'h918)
`define CLP_KV_REG_KEY_ENTRY_16_7                                                                   (32'h1001891c)
`define KV_REG_KEY_ENTRY_16_7                                                                       (32'h91c)
`define CLP_KV_REG_KEY_ENTRY_16_8                                                                   (32'h10018920)
`define KV_REG_KEY_ENTRY_16_8                                                                       (32'h920)
`define CLP_KV_REG_KEY_ENTRY_16_9                                                                   (32'h10018924)
`define KV_REG_KEY_ENTRY_16_9                                                                       (32'h924)
`define CLP_KV_REG_KEY_ENTRY_16_10                                                                  (32'h10018928)
`define KV_REG_KEY_ENTRY_16_10                                                                      (32'h928)
`define CLP_KV_REG_KEY_ENTRY_16_11                                                                  (32'h1001892c)
`define KV_REG_KEY_ENTRY_16_11                                                                      (32'h92c)
`define CLP_KV_REG_KEY_ENTRY_17_0                                                                   (32'h10018930)
`define KV_REG_KEY_ENTRY_17_0                                                                       (32'h930)
`define CLP_KV_REG_KEY_ENTRY_17_1                                                                   (32'h10018934)
`define KV_REG_KEY_ENTRY_17_1                                                                       (32'h934)
`define CLP_KV_REG_KEY_ENTRY_17_2                                                                   (32'h10018938)
`define KV_REG_KEY_ENTRY_17_2                                                                       (32'h938)
`define CLP_KV_REG_KEY_ENTRY_17_3                                                                   (32'h1001893c)
`define KV_REG_KEY_ENTRY_17_3                                                                       (32'h93c)
`define CLP_KV_REG_KEY_ENTRY_17_4                                                                   (32'h10018940)
`define KV_REG_KEY_ENTRY_17_4                                                                       (32'h940)
`define CLP_KV_REG_KEY_ENTRY_17_5                                                                   (32'h10018944)
`define KV_REG_KEY_ENTRY_17_5                                                                       (32'h944)
`define CLP_KV_REG_KEY_ENTRY_17_6                                                                   (32'h10018948)
`define KV_REG_KEY_ENTRY_17_6                                                                       (32'h948)
`define CLP_KV_REG_KEY_ENTRY_17_7                                                                   (32'h1001894c)
`define KV_REG_KEY_ENTRY_17_7                                                                       (32'h94c)
`define CLP_KV_REG_KEY_ENTRY_17_8                                                                   (32'h10018950)
`define KV_REG_KEY_ENTRY_17_8                                                                       (32'h950)
`define CLP_KV_REG_KEY_ENTRY_17_9                                                                   (32'h10018954)
`define KV_REG_KEY_ENTRY_17_9                                                                       (32'h954)
`define CLP_KV_REG_KEY_ENTRY_17_10                                                                  (32'h10018958)
`define KV_REG_KEY_ENTRY_17_10                                                                      (32'h958)
`define CLP_KV_REG_KEY_ENTRY_17_11                                                                  (32'h1001895c)
`define KV_REG_KEY_ENTRY_17_11                                                                      (32'h95c)
`define CLP_KV_REG_KEY_ENTRY_18_0                                                                   (32'h10018960)
`define KV_REG_KEY_ENTRY_18_0                                                                       (32'h960)
`define CLP_KV_REG_KEY_ENTRY_18_1                                                                   (32'h10018964)
`define KV_REG_KEY_ENTRY_18_1                                                                       (32'h964)
`define CLP_KV_REG_KEY_ENTRY_18_2                                                                   (32'h10018968)
`define KV_REG_KEY_ENTRY_18_2                                                                       (32'h968)
`define CLP_KV_REG_KEY_ENTRY_18_3                                                                   (32'h1001896c)
`define KV_REG_KEY_ENTRY_18_3                                                                       (32'h96c)
`define CLP_KV_REG_KEY_ENTRY_18_4                                                                   (32'h10018970)
`define KV_REG_KEY_ENTRY_18_4                                                                       (32'h970)
`define CLP_KV_REG_KEY_ENTRY_18_5                                                                   (32'h10018974)
`define KV_REG_KEY_ENTRY_18_5                                                                       (32'h974)
`define CLP_KV_REG_KEY_ENTRY_18_6                                                                   (32'h10018978)
`define KV_REG_KEY_ENTRY_18_6                                                                       (32'h978)
`define CLP_KV_REG_KEY_ENTRY_18_7                                                                   (32'h1001897c)
`define KV_REG_KEY_ENTRY_18_7                                                                       (32'h97c)
`define CLP_KV_REG_KEY_ENTRY_18_8                                                                   (32'h10018980)
`define KV_REG_KEY_ENTRY_18_8                                                                       (32'h980)
`define CLP_KV_REG_KEY_ENTRY_18_9                                                                   (32'h10018984)
`define KV_REG_KEY_ENTRY_18_9                                                                       (32'h984)
`define CLP_KV_REG_KEY_ENTRY_18_10                                                                  (32'h10018988)
`define KV_REG_KEY_ENTRY_18_10                                                                      (32'h988)
`define CLP_KV_REG_KEY_ENTRY_18_11                                                                  (32'h1001898c)
`define KV_REG_KEY_ENTRY_18_11                                                                      (32'h98c)
`define CLP_KV_REG_KEY_ENTRY_19_0                                                                   (32'h10018990)
`define KV_REG_KEY_ENTRY_19_0                                                                       (32'h990)
`define CLP_KV_REG_KEY_ENTRY_19_1                                                                   (32'h10018994)
`define KV_REG_KEY_ENTRY_19_1                                                                       (32'h994)
`define CLP_KV_REG_KEY_ENTRY_19_2                                                                   (32'h10018998)
`define KV_REG_KEY_ENTRY_19_2                                                                       (32'h998)
`define CLP_KV_REG_KEY_ENTRY_19_3                                                                   (32'h1001899c)
`define KV_REG_KEY_ENTRY_19_3                                                                       (32'h99c)
`define CLP_KV_REG_KEY_ENTRY_19_4                                                                   (32'h100189a0)
`define KV_REG_KEY_ENTRY_19_4                                                                       (32'h9a0)
`define CLP_KV_REG_KEY_ENTRY_19_5                                                                   (32'h100189a4)
`define KV_REG_KEY_ENTRY_19_5                                                                       (32'h9a4)
`define CLP_KV_REG_KEY_ENTRY_19_6                                                                   (32'h100189a8)
`define KV_REG_KEY_ENTRY_19_6                                                                       (32'h9a8)
`define CLP_KV_REG_KEY_ENTRY_19_7                                                                   (32'h100189ac)
`define KV_REG_KEY_ENTRY_19_7                                                                       (32'h9ac)
`define CLP_KV_REG_KEY_ENTRY_19_8                                                                   (32'h100189b0)
`define KV_REG_KEY_ENTRY_19_8                                                                       (32'h9b0)
`define CLP_KV_REG_KEY_ENTRY_19_9                                                                   (32'h100189b4)
`define KV_REG_KEY_ENTRY_19_9                                                                       (32'h9b4)
`define CLP_KV_REG_KEY_ENTRY_19_10                                                                  (32'h100189b8)
`define KV_REG_KEY_ENTRY_19_10                                                                      (32'h9b8)
`define CLP_KV_REG_KEY_ENTRY_19_11                                                                  (32'h100189bc)
`define KV_REG_KEY_ENTRY_19_11                                                                      (32'h9bc)
`define CLP_KV_REG_KEY_ENTRY_20_0                                                                   (32'h100189c0)
`define KV_REG_KEY_ENTRY_20_0                                                                       (32'h9c0)
`define CLP_KV_REG_KEY_ENTRY_20_1                                                                   (32'h100189c4)
`define KV_REG_KEY_ENTRY_20_1                                                                       (32'h9c4)
`define CLP_KV_REG_KEY_ENTRY_20_2                                                                   (32'h100189c8)
`define KV_REG_KEY_ENTRY_20_2                                                                       (32'h9c8)
`define CLP_KV_REG_KEY_ENTRY_20_3                                                                   (32'h100189cc)
`define KV_REG_KEY_ENTRY_20_3                                                                       (32'h9cc)
`define CLP_KV_REG_KEY_ENTRY_20_4                                                                   (32'h100189d0)
`define KV_REG_KEY_ENTRY_20_4                                                                       (32'h9d0)
`define CLP_KV_REG_KEY_ENTRY_20_5                                                                   (32'h100189d4)
`define KV_REG_KEY_ENTRY_20_5                                                                       (32'h9d4)
`define CLP_KV_REG_KEY_ENTRY_20_6                                                                   (32'h100189d8)
`define KV_REG_KEY_ENTRY_20_6                                                                       (32'h9d8)
`define CLP_KV_REG_KEY_ENTRY_20_7                                                                   (32'h100189dc)
`define KV_REG_KEY_ENTRY_20_7                                                                       (32'h9dc)
`define CLP_KV_REG_KEY_ENTRY_20_8                                                                   (32'h100189e0)
`define KV_REG_KEY_ENTRY_20_8                                                                       (32'h9e0)
`define CLP_KV_REG_KEY_ENTRY_20_9                                                                   (32'h100189e4)
`define KV_REG_KEY_ENTRY_20_9                                                                       (32'h9e4)
`define CLP_KV_REG_KEY_ENTRY_20_10                                                                  (32'h100189e8)
`define KV_REG_KEY_ENTRY_20_10                                                                      (32'h9e8)
`define CLP_KV_REG_KEY_ENTRY_20_11                                                                  (32'h100189ec)
`define KV_REG_KEY_ENTRY_20_11                                                                      (32'h9ec)
`define CLP_KV_REG_KEY_ENTRY_21_0                                                                   (32'h100189f0)
`define KV_REG_KEY_ENTRY_21_0                                                                       (32'h9f0)
`define CLP_KV_REG_KEY_ENTRY_21_1                                                                   (32'h100189f4)
`define KV_REG_KEY_ENTRY_21_1                                                                       (32'h9f4)
`define CLP_KV_REG_KEY_ENTRY_21_2                                                                   (32'h100189f8)
`define KV_REG_KEY_ENTRY_21_2                                                                       (32'h9f8)
`define CLP_KV_REG_KEY_ENTRY_21_3                                                                   (32'h100189fc)
`define KV_REG_KEY_ENTRY_21_3                                                                       (32'h9fc)
`define CLP_KV_REG_KEY_ENTRY_21_4                                                                   (32'h10018a00)
`define KV_REG_KEY_ENTRY_21_4                                                                       (32'ha00)
`define CLP_KV_REG_KEY_ENTRY_21_5                                                                   (32'h10018a04)
`define KV_REG_KEY_ENTRY_21_5                                                                       (32'ha04)
`define CLP_KV_REG_KEY_ENTRY_21_6                                                                   (32'h10018a08)
`define KV_REG_KEY_ENTRY_21_6                                                                       (32'ha08)
`define CLP_KV_REG_KEY_ENTRY_21_7                                                                   (32'h10018a0c)
`define KV_REG_KEY_ENTRY_21_7                                                                       (32'ha0c)
`define CLP_KV_REG_KEY_ENTRY_21_8                                                                   (32'h10018a10)
`define KV_REG_KEY_ENTRY_21_8                                                                       (32'ha10)
`define CLP_KV_REG_KEY_ENTRY_21_9                                                                   (32'h10018a14)
`define KV_REG_KEY_ENTRY_21_9                                                                       (32'ha14)
`define CLP_KV_REG_KEY_ENTRY_21_10                                                                  (32'h10018a18)
`define KV_REG_KEY_ENTRY_21_10                                                                      (32'ha18)
`define CLP_KV_REG_KEY_ENTRY_21_11                                                                  (32'h10018a1c)
`define KV_REG_KEY_ENTRY_21_11                                                                      (32'ha1c)
`define CLP_KV_REG_KEY_ENTRY_22_0                                                                   (32'h10018a20)
`define KV_REG_KEY_ENTRY_22_0                                                                       (32'ha20)
`define CLP_KV_REG_KEY_ENTRY_22_1                                                                   (32'h10018a24)
`define KV_REG_KEY_ENTRY_22_1                                                                       (32'ha24)
`define CLP_KV_REG_KEY_ENTRY_22_2                                                                   (32'h10018a28)
`define KV_REG_KEY_ENTRY_22_2                                                                       (32'ha28)
`define CLP_KV_REG_KEY_ENTRY_22_3                                                                   (32'h10018a2c)
`define KV_REG_KEY_ENTRY_22_3                                                                       (32'ha2c)
`define CLP_KV_REG_KEY_ENTRY_22_4                                                                   (32'h10018a30)
`define KV_REG_KEY_ENTRY_22_4                                                                       (32'ha30)
`define CLP_KV_REG_KEY_ENTRY_22_5                                                                   (32'h10018a34)
`define KV_REG_KEY_ENTRY_22_5                                                                       (32'ha34)
`define CLP_KV_REG_KEY_ENTRY_22_6                                                                   (32'h10018a38)
`define KV_REG_KEY_ENTRY_22_6                                                                       (32'ha38)
`define CLP_KV_REG_KEY_ENTRY_22_7                                                                   (32'h10018a3c)
`define KV_REG_KEY_ENTRY_22_7                                                                       (32'ha3c)
`define CLP_KV_REG_KEY_ENTRY_22_8                                                                   (32'h10018a40)
`define KV_REG_KEY_ENTRY_22_8                                                                       (32'ha40)
`define CLP_KV_REG_KEY_ENTRY_22_9                                                                   (32'h10018a44)
`define KV_REG_KEY_ENTRY_22_9                                                                       (32'ha44)
`define CLP_KV_REG_KEY_ENTRY_22_10                                                                  (32'h10018a48)
`define KV_REG_KEY_ENTRY_22_10                                                                      (32'ha48)
`define CLP_KV_REG_KEY_ENTRY_22_11                                                                  (32'h10018a4c)
`define KV_REG_KEY_ENTRY_22_11                                                                      (32'ha4c)
`define CLP_KV_REG_KEY_ENTRY_23_0                                                                   (32'h10018a50)
`define KV_REG_KEY_ENTRY_23_0                                                                       (32'ha50)
`define CLP_KV_REG_KEY_ENTRY_23_1                                                                   (32'h10018a54)
`define KV_REG_KEY_ENTRY_23_1                                                                       (32'ha54)
`define CLP_KV_REG_KEY_ENTRY_23_2                                                                   (32'h10018a58)
`define KV_REG_KEY_ENTRY_23_2                                                                       (32'ha58)
`define CLP_KV_REG_KEY_ENTRY_23_3                                                                   (32'h10018a5c)
`define KV_REG_KEY_ENTRY_23_3                                                                       (32'ha5c)
`define CLP_KV_REG_KEY_ENTRY_23_4                                                                   (32'h10018a60)
`define KV_REG_KEY_ENTRY_23_4                                                                       (32'ha60)
`define CLP_KV_REG_KEY_ENTRY_23_5                                                                   (32'h10018a64)
`define KV_REG_KEY_ENTRY_23_5                                                                       (32'ha64)
`define CLP_KV_REG_KEY_ENTRY_23_6                                                                   (32'h10018a68)
`define KV_REG_KEY_ENTRY_23_6                                                                       (32'ha68)
`define CLP_KV_REG_KEY_ENTRY_23_7                                                                   (32'h10018a6c)
`define KV_REG_KEY_ENTRY_23_7                                                                       (32'ha6c)
`define CLP_KV_REG_KEY_ENTRY_23_8                                                                   (32'h10018a70)
`define KV_REG_KEY_ENTRY_23_8                                                                       (32'ha70)
`define CLP_KV_REG_KEY_ENTRY_23_9                                                                   (32'h10018a74)
`define KV_REG_KEY_ENTRY_23_9                                                                       (32'ha74)
`define CLP_KV_REG_KEY_ENTRY_23_10                                                                  (32'h10018a78)
`define KV_REG_KEY_ENTRY_23_10                                                                      (32'ha78)
`define CLP_KV_REG_KEY_ENTRY_23_11                                                                  (32'h10018a7c)
`define KV_REG_KEY_ENTRY_23_11                                                                      (32'ha7c)
`define CLP_KV_REG_KEY_ENTRY_24_0                                                                   (32'h10018a80)
`define KV_REG_KEY_ENTRY_24_0                                                                       (32'ha80)
`define CLP_KV_REG_KEY_ENTRY_24_1                                                                   (32'h10018a84)
`define KV_REG_KEY_ENTRY_24_1                                                                       (32'ha84)
`define CLP_KV_REG_KEY_ENTRY_24_2                                                                   (32'h10018a88)
`define KV_REG_KEY_ENTRY_24_2                                                                       (32'ha88)
`define CLP_KV_REG_KEY_ENTRY_24_3                                                                   (32'h10018a8c)
`define KV_REG_KEY_ENTRY_24_3                                                                       (32'ha8c)
`define CLP_KV_REG_KEY_ENTRY_24_4                                                                   (32'h10018a90)
`define KV_REG_KEY_ENTRY_24_4                                                                       (32'ha90)
`define CLP_KV_REG_KEY_ENTRY_24_5                                                                   (32'h10018a94)
`define KV_REG_KEY_ENTRY_24_5                                                                       (32'ha94)
`define CLP_KV_REG_KEY_ENTRY_24_6                                                                   (32'h10018a98)
`define KV_REG_KEY_ENTRY_24_6                                                                       (32'ha98)
`define CLP_KV_REG_KEY_ENTRY_24_7                                                                   (32'h10018a9c)
`define KV_REG_KEY_ENTRY_24_7                                                                       (32'ha9c)
`define CLP_KV_REG_KEY_ENTRY_24_8                                                                   (32'h10018aa0)
`define KV_REG_KEY_ENTRY_24_8                                                                       (32'haa0)
`define CLP_KV_REG_KEY_ENTRY_24_9                                                                   (32'h10018aa4)
`define KV_REG_KEY_ENTRY_24_9                                                                       (32'haa4)
`define CLP_KV_REG_KEY_ENTRY_24_10                                                                  (32'h10018aa8)
`define KV_REG_KEY_ENTRY_24_10                                                                      (32'haa8)
`define CLP_KV_REG_KEY_ENTRY_24_11                                                                  (32'h10018aac)
`define KV_REG_KEY_ENTRY_24_11                                                                      (32'haac)
`define CLP_KV_REG_KEY_ENTRY_25_0                                                                   (32'h10018ab0)
`define KV_REG_KEY_ENTRY_25_0                                                                       (32'hab0)
`define CLP_KV_REG_KEY_ENTRY_25_1                                                                   (32'h10018ab4)
`define KV_REG_KEY_ENTRY_25_1                                                                       (32'hab4)
`define CLP_KV_REG_KEY_ENTRY_25_2                                                                   (32'h10018ab8)
`define KV_REG_KEY_ENTRY_25_2                                                                       (32'hab8)
`define CLP_KV_REG_KEY_ENTRY_25_3                                                                   (32'h10018abc)
`define KV_REG_KEY_ENTRY_25_3                                                                       (32'habc)
`define CLP_KV_REG_KEY_ENTRY_25_4                                                                   (32'h10018ac0)
`define KV_REG_KEY_ENTRY_25_4                                                                       (32'hac0)
`define CLP_KV_REG_KEY_ENTRY_25_5                                                                   (32'h10018ac4)
`define KV_REG_KEY_ENTRY_25_5                                                                       (32'hac4)
`define CLP_KV_REG_KEY_ENTRY_25_6                                                                   (32'h10018ac8)
`define KV_REG_KEY_ENTRY_25_6                                                                       (32'hac8)
`define CLP_KV_REG_KEY_ENTRY_25_7                                                                   (32'h10018acc)
`define KV_REG_KEY_ENTRY_25_7                                                                       (32'hacc)
`define CLP_KV_REG_KEY_ENTRY_25_8                                                                   (32'h10018ad0)
`define KV_REG_KEY_ENTRY_25_8                                                                       (32'had0)
`define CLP_KV_REG_KEY_ENTRY_25_9                                                                   (32'h10018ad4)
`define KV_REG_KEY_ENTRY_25_9                                                                       (32'had4)
`define CLP_KV_REG_KEY_ENTRY_25_10                                                                  (32'h10018ad8)
`define KV_REG_KEY_ENTRY_25_10                                                                      (32'had8)
`define CLP_KV_REG_KEY_ENTRY_25_11                                                                  (32'h10018adc)
`define KV_REG_KEY_ENTRY_25_11                                                                      (32'hadc)
`define CLP_KV_REG_KEY_ENTRY_26_0                                                                   (32'h10018ae0)
`define KV_REG_KEY_ENTRY_26_0                                                                       (32'hae0)
`define CLP_KV_REG_KEY_ENTRY_26_1                                                                   (32'h10018ae4)
`define KV_REG_KEY_ENTRY_26_1                                                                       (32'hae4)
`define CLP_KV_REG_KEY_ENTRY_26_2                                                                   (32'h10018ae8)
`define KV_REG_KEY_ENTRY_26_2                                                                       (32'hae8)
`define CLP_KV_REG_KEY_ENTRY_26_3                                                                   (32'h10018aec)
`define KV_REG_KEY_ENTRY_26_3                                                                       (32'haec)
`define CLP_KV_REG_KEY_ENTRY_26_4                                                                   (32'h10018af0)
`define KV_REG_KEY_ENTRY_26_4                                                                       (32'haf0)
`define CLP_KV_REG_KEY_ENTRY_26_5                                                                   (32'h10018af4)
`define KV_REG_KEY_ENTRY_26_5                                                                       (32'haf4)
`define CLP_KV_REG_KEY_ENTRY_26_6                                                                   (32'h10018af8)
`define KV_REG_KEY_ENTRY_26_6                                                                       (32'haf8)
`define CLP_KV_REG_KEY_ENTRY_26_7                                                                   (32'h10018afc)
`define KV_REG_KEY_ENTRY_26_7                                                                       (32'hafc)
`define CLP_KV_REG_KEY_ENTRY_26_8                                                                   (32'h10018b00)
`define KV_REG_KEY_ENTRY_26_8                                                                       (32'hb00)
`define CLP_KV_REG_KEY_ENTRY_26_9                                                                   (32'h10018b04)
`define KV_REG_KEY_ENTRY_26_9                                                                       (32'hb04)
`define CLP_KV_REG_KEY_ENTRY_26_10                                                                  (32'h10018b08)
`define KV_REG_KEY_ENTRY_26_10                                                                      (32'hb08)
`define CLP_KV_REG_KEY_ENTRY_26_11                                                                  (32'h10018b0c)
`define KV_REG_KEY_ENTRY_26_11                                                                      (32'hb0c)
`define CLP_KV_REG_KEY_ENTRY_27_0                                                                   (32'h10018b10)
`define KV_REG_KEY_ENTRY_27_0                                                                       (32'hb10)
`define CLP_KV_REG_KEY_ENTRY_27_1                                                                   (32'h10018b14)
`define KV_REG_KEY_ENTRY_27_1                                                                       (32'hb14)
`define CLP_KV_REG_KEY_ENTRY_27_2                                                                   (32'h10018b18)
`define KV_REG_KEY_ENTRY_27_2                                                                       (32'hb18)
`define CLP_KV_REG_KEY_ENTRY_27_3                                                                   (32'h10018b1c)
`define KV_REG_KEY_ENTRY_27_3                                                                       (32'hb1c)
`define CLP_KV_REG_KEY_ENTRY_27_4                                                                   (32'h10018b20)
`define KV_REG_KEY_ENTRY_27_4                                                                       (32'hb20)
`define CLP_KV_REG_KEY_ENTRY_27_5                                                                   (32'h10018b24)
`define KV_REG_KEY_ENTRY_27_5                                                                       (32'hb24)
`define CLP_KV_REG_KEY_ENTRY_27_6                                                                   (32'h10018b28)
`define KV_REG_KEY_ENTRY_27_6                                                                       (32'hb28)
`define CLP_KV_REG_KEY_ENTRY_27_7                                                                   (32'h10018b2c)
`define KV_REG_KEY_ENTRY_27_7                                                                       (32'hb2c)
`define CLP_KV_REG_KEY_ENTRY_27_8                                                                   (32'h10018b30)
`define KV_REG_KEY_ENTRY_27_8                                                                       (32'hb30)
`define CLP_KV_REG_KEY_ENTRY_27_9                                                                   (32'h10018b34)
`define KV_REG_KEY_ENTRY_27_9                                                                       (32'hb34)
`define CLP_KV_REG_KEY_ENTRY_27_10                                                                  (32'h10018b38)
`define KV_REG_KEY_ENTRY_27_10                                                                      (32'hb38)
`define CLP_KV_REG_KEY_ENTRY_27_11                                                                  (32'h10018b3c)
`define KV_REG_KEY_ENTRY_27_11                                                                      (32'hb3c)
`define CLP_KV_REG_KEY_ENTRY_28_0                                                                   (32'h10018b40)
`define KV_REG_KEY_ENTRY_28_0                                                                       (32'hb40)
`define CLP_KV_REG_KEY_ENTRY_28_1                                                                   (32'h10018b44)
`define KV_REG_KEY_ENTRY_28_1                                                                       (32'hb44)
`define CLP_KV_REG_KEY_ENTRY_28_2                                                                   (32'h10018b48)
`define KV_REG_KEY_ENTRY_28_2                                                                       (32'hb48)
`define CLP_KV_REG_KEY_ENTRY_28_3                                                                   (32'h10018b4c)
`define KV_REG_KEY_ENTRY_28_3                                                                       (32'hb4c)
`define CLP_KV_REG_KEY_ENTRY_28_4                                                                   (32'h10018b50)
`define KV_REG_KEY_ENTRY_28_4                                                                       (32'hb50)
`define CLP_KV_REG_KEY_ENTRY_28_5                                                                   (32'h10018b54)
`define KV_REG_KEY_ENTRY_28_5                                                                       (32'hb54)
`define CLP_KV_REG_KEY_ENTRY_28_6                                                                   (32'h10018b58)
`define KV_REG_KEY_ENTRY_28_6                                                                       (32'hb58)
`define CLP_KV_REG_KEY_ENTRY_28_7                                                                   (32'h10018b5c)
`define KV_REG_KEY_ENTRY_28_7                                                                       (32'hb5c)
`define CLP_KV_REG_KEY_ENTRY_28_8                                                                   (32'h10018b60)
`define KV_REG_KEY_ENTRY_28_8                                                                       (32'hb60)
`define CLP_KV_REG_KEY_ENTRY_28_9                                                                   (32'h10018b64)
`define KV_REG_KEY_ENTRY_28_9                                                                       (32'hb64)
`define CLP_KV_REG_KEY_ENTRY_28_10                                                                  (32'h10018b68)
`define KV_REG_KEY_ENTRY_28_10                                                                      (32'hb68)
`define CLP_KV_REG_KEY_ENTRY_28_11                                                                  (32'h10018b6c)
`define KV_REG_KEY_ENTRY_28_11                                                                      (32'hb6c)
`define CLP_KV_REG_KEY_ENTRY_29_0                                                                   (32'h10018b70)
`define KV_REG_KEY_ENTRY_29_0                                                                       (32'hb70)
`define CLP_KV_REG_KEY_ENTRY_29_1                                                                   (32'h10018b74)
`define KV_REG_KEY_ENTRY_29_1                                                                       (32'hb74)
`define CLP_KV_REG_KEY_ENTRY_29_2                                                                   (32'h10018b78)
`define KV_REG_KEY_ENTRY_29_2                                                                       (32'hb78)
`define CLP_KV_REG_KEY_ENTRY_29_3                                                                   (32'h10018b7c)
`define KV_REG_KEY_ENTRY_29_3                                                                       (32'hb7c)
`define CLP_KV_REG_KEY_ENTRY_29_4                                                                   (32'h10018b80)
`define KV_REG_KEY_ENTRY_29_4                                                                       (32'hb80)
`define CLP_KV_REG_KEY_ENTRY_29_5                                                                   (32'h10018b84)
`define KV_REG_KEY_ENTRY_29_5                                                                       (32'hb84)
`define CLP_KV_REG_KEY_ENTRY_29_6                                                                   (32'h10018b88)
`define KV_REG_KEY_ENTRY_29_6                                                                       (32'hb88)
`define CLP_KV_REG_KEY_ENTRY_29_7                                                                   (32'h10018b8c)
`define KV_REG_KEY_ENTRY_29_7                                                                       (32'hb8c)
`define CLP_KV_REG_KEY_ENTRY_29_8                                                                   (32'h10018b90)
`define KV_REG_KEY_ENTRY_29_8                                                                       (32'hb90)
`define CLP_KV_REG_KEY_ENTRY_29_9                                                                   (32'h10018b94)
`define KV_REG_KEY_ENTRY_29_9                                                                       (32'hb94)
`define CLP_KV_REG_KEY_ENTRY_29_10                                                                  (32'h10018b98)
`define KV_REG_KEY_ENTRY_29_10                                                                      (32'hb98)
`define CLP_KV_REG_KEY_ENTRY_29_11                                                                  (32'h10018b9c)
`define KV_REG_KEY_ENTRY_29_11                                                                      (32'hb9c)
`define CLP_KV_REG_KEY_ENTRY_30_0                                                                   (32'h10018ba0)
`define KV_REG_KEY_ENTRY_30_0                                                                       (32'hba0)
`define CLP_KV_REG_KEY_ENTRY_30_1                                                                   (32'h10018ba4)
`define KV_REG_KEY_ENTRY_30_1                                                                       (32'hba4)
`define CLP_KV_REG_KEY_ENTRY_30_2                                                                   (32'h10018ba8)
`define KV_REG_KEY_ENTRY_30_2                                                                       (32'hba8)
`define CLP_KV_REG_KEY_ENTRY_30_3                                                                   (32'h10018bac)
`define KV_REG_KEY_ENTRY_30_3                                                                       (32'hbac)
`define CLP_KV_REG_KEY_ENTRY_30_4                                                                   (32'h10018bb0)
`define KV_REG_KEY_ENTRY_30_4                                                                       (32'hbb0)
`define CLP_KV_REG_KEY_ENTRY_30_5                                                                   (32'h10018bb4)
`define KV_REG_KEY_ENTRY_30_5                                                                       (32'hbb4)
`define CLP_KV_REG_KEY_ENTRY_30_6                                                                   (32'h10018bb8)
`define KV_REG_KEY_ENTRY_30_6                                                                       (32'hbb8)
`define CLP_KV_REG_KEY_ENTRY_30_7                                                                   (32'h10018bbc)
`define KV_REG_KEY_ENTRY_30_7                                                                       (32'hbbc)
`define CLP_KV_REG_KEY_ENTRY_30_8                                                                   (32'h10018bc0)
`define KV_REG_KEY_ENTRY_30_8                                                                       (32'hbc0)
`define CLP_KV_REG_KEY_ENTRY_30_9                                                                   (32'h10018bc4)
`define KV_REG_KEY_ENTRY_30_9                                                                       (32'hbc4)
`define CLP_KV_REG_KEY_ENTRY_30_10                                                                  (32'h10018bc8)
`define KV_REG_KEY_ENTRY_30_10                                                                      (32'hbc8)
`define CLP_KV_REG_KEY_ENTRY_30_11                                                                  (32'h10018bcc)
`define KV_REG_KEY_ENTRY_30_11                                                                      (32'hbcc)
`define CLP_KV_REG_KEY_ENTRY_31_0                                                                   (32'h10018bd0)
`define KV_REG_KEY_ENTRY_31_0                                                                       (32'hbd0)
`define CLP_KV_REG_KEY_ENTRY_31_1                                                                   (32'h10018bd4)
`define KV_REG_KEY_ENTRY_31_1                                                                       (32'hbd4)
`define CLP_KV_REG_KEY_ENTRY_31_2                                                                   (32'h10018bd8)
`define KV_REG_KEY_ENTRY_31_2                                                                       (32'hbd8)
`define CLP_KV_REG_KEY_ENTRY_31_3                                                                   (32'h10018bdc)
`define KV_REG_KEY_ENTRY_31_3                                                                       (32'hbdc)
`define CLP_KV_REG_KEY_ENTRY_31_4                                                                   (32'h10018be0)
`define KV_REG_KEY_ENTRY_31_4                                                                       (32'hbe0)
`define CLP_KV_REG_KEY_ENTRY_31_5                                                                   (32'h10018be4)
`define KV_REG_KEY_ENTRY_31_5                                                                       (32'hbe4)
`define CLP_KV_REG_KEY_ENTRY_31_6                                                                   (32'h10018be8)
`define KV_REG_KEY_ENTRY_31_6                                                                       (32'hbe8)
`define CLP_KV_REG_KEY_ENTRY_31_7                                                                   (32'h10018bec)
`define KV_REG_KEY_ENTRY_31_7                                                                       (32'hbec)
`define CLP_KV_REG_KEY_ENTRY_31_8                                                                   (32'h10018bf0)
`define KV_REG_KEY_ENTRY_31_8                                                                       (32'hbf0)
`define CLP_KV_REG_KEY_ENTRY_31_9                                                                   (32'h10018bf4)
`define KV_REG_KEY_ENTRY_31_9                                                                       (32'hbf4)
`define CLP_KV_REG_KEY_ENTRY_31_10                                                                  (32'h10018bf8)
`define KV_REG_KEY_ENTRY_31_10                                                                      (32'hbf8)
`define CLP_KV_REG_KEY_ENTRY_31_11                                                                  (32'h10018bfc)
`define KV_REG_KEY_ENTRY_31_11                                                                      (32'hbfc)
`define CLP_KV_REG_CLEAR_SECRETS                                                                    (32'h10018c00)
`define KV_REG_CLEAR_SECRETS                                                                        (32'hc00)
`define KV_REG_CLEAR_SECRETS_WR_DEBUG_VALUES_LOW                                                    (0)
`define KV_REG_CLEAR_SECRETS_WR_DEBUG_VALUES_MASK                                                   (32'h1)
`define KV_REG_CLEAR_SECRETS_SEL_DEBUG_VALUE_LOW                                                    (1)
`define KV_REG_CLEAR_SECRETS_SEL_DEBUG_VALUE_MASK                                                   (32'h2)
`define CLP_PV_REG_BASE_ADDR                                                                        (32'h1001a000)
`define CLP_PV_REG_PCR_CTRL_0                                                                       (32'h1001a000)
`define PV_REG_PCR_CTRL_0                                                                           (32'h0)
`define PV_REG_PCR_CTRL_0_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_0_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_0_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_0_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_0_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_0_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_0_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_0_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_1                                                                       (32'h1001a004)
`define PV_REG_PCR_CTRL_1                                                                           (32'h4)
`define PV_REG_PCR_CTRL_1_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_1_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_1_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_1_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_1_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_1_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_1_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_1_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_2                                                                       (32'h1001a008)
`define PV_REG_PCR_CTRL_2                                                                           (32'h8)
`define PV_REG_PCR_CTRL_2_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_2_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_2_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_2_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_2_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_2_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_2_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_2_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_3                                                                       (32'h1001a00c)
`define PV_REG_PCR_CTRL_3                                                                           (32'hc)
`define PV_REG_PCR_CTRL_3_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_3_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_3_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_3_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_3_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_3_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_3_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_3_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_4                                                                       (32'h1001a010)
`define PV_REG_PCR_CTRL_4                                                                           (32'h10)
`define PV_REG_PCR_CTRL_4_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_4_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_4_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_4_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_4_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_4_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_4_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_4_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_5                                                                       (32'h1001a014)
`define PV_REG_PCR_CTRL_5                                                                           (32'h14)
`define PV_REG_PCR_CTRL_5_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_5_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_5_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_5_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_5_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_5_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_5_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_5_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_6                                                                       (32'h1001a018)
`define PV_REG_PCR_CTRL_6                                                                           (32'h18)
`define PV_REG_PCR_CTRL_6_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_6_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_6_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_6_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_6_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_6_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_6_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_6_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_7                                                                       (32'h1001a01c)
`define PV_REG_PCR_CTRL_7                                                                           (32'h1c)
`define PV_REG_PCR_CTRL_7_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_7_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_7_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_7_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_7_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_7_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_7_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_7_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_8                                                                       (32'h1001a020)
`define PV_REG_PCR_CTRL_8                                                                           (32'h20)
`define PV_REG_PCR_CTRL_8_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_8_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_8_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_8_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_8_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_8_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_8_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_8_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_9                                                                       (32'h1001a024)
`define PV_REG_PCR_CTRL_9                                                                           (32'h24)
`define PV_REG_PCR_CTRL_9_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_9_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_9_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_9_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_9_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_9_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_9_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_9_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_10                                                                      (32'h1001a028)
`define PV_REG_PCR_CTRL_10                                                                          (32'h28)
`define PV_REG_PCR_CTRL_10_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_10_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_10_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_10_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_10_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_10_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_10_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_10_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_11                                                                      (32'h1001a02c)
`define PV_REG_PCR_CTRL_11                                                                          (32'h2c)
`define PV_REG_PCR_CTRL_11_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_11_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_11_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_11_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_11_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_11_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_11_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_11_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_12                                                                      (32'h1001a030)
`define PV_REG_PCR_CTRL_12                                                                          (32'h30)
`define PV_REG_PCR_CTRL_12_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_12_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_12_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_12_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_12_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_12_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_12_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_12_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_13                                                                      (32'h1001a034)
`define PV_REG_PCR_CTRL_13                                                                          (32'h34)
`define PV_REG_PCR_CTRL_13_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_13_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_13_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_13_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_13_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_13_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_13_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_13_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_14                                                                      (32'h1001a038)
`define PV_REG_PCR_CTRL_14                                                                          (32'h38)
`define PV_REG_PCR_CTRL_14_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_14_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_14_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_14_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_14_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_14_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_14_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_14_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_15                                                                      (32'h1001a03c)
`define PV_REG_PCR_CTRL_15                                                                          (32'h3c)
`define PV_REG_PCR_CTRL_15_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_15_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_15_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_15_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_15_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_15_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_15_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_15_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_16                                                                      (32'h1001a040)
`define PV_REG_PCR_CTRL_16                                                                          (32'h40)
`define PV_REG_PCR_CTRL_16_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_16_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_16_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_16_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_16_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_16_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_16_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_16_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_17                                                                      (32'h1001a044)
`define PV_REG_PCR_CTRL_17                                                                          (32'h44)
`define PV_REG_PCR_CTRL_17_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_17_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_17_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_17_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_17_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_17_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_17_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_17_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_18                                                                      (32'h1001a048)
`define PV_REG_PCR_CTRL_18                                                                          (32'h48)
`define PV_REG_PCR_CTRL_18_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_18_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_18_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_18_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_18_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_18_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_18_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_18_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_19                                                                      (32'h1001a04c)
`define PV_REG_PCR_CTRL_19                                                                          (32'h4c)
`define PV_REG_PCR_CTRL_19_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_19_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_19_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_19_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_19_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_19_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_19_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_19_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_20                                                                      (32'h1001a050)
`define PV_REG_PCR_CTRL_20                                                                          (32'h50)
`define PV_REG_PCR_CTRL_20_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_20_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_20_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_20_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_20_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_20_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_20_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_20_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_21                                                                      (32'h1001a054)
`define PV_REG_PCR_CTRL_21                                                                          (32'h54)
`define PV_REG_PCR_CTRL_21_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_21_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_21_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_21_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_21_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_21_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_21_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_21_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_22                                                                      (32'h1001a058)
`define PV_REG_PCR_CTRL_22                                                                          (32'h58)
`define PV_REG_PCR_CTRL_22_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_22_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_22_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_22_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_22_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_22_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_22_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_22_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_23                                                                      (32'h1001a05c)
`define PV_REG_PCR_CTRL_23                                                                          (32'h5c)
`define PV_REG_PCR_CTRL_23_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_23_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_23_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_23_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_23_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_23_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_23_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_23_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_24                                                                      (32'h1001a060)
`define PV_REG_PCR_CTRL_24                                                                          (32'h60)
`define PV_REG_PCR_CTRL_24_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_24_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_24_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_24_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_24_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_24_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_24_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_24_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_25                                                                      (32'h1001a064)
`define PV_REG_PCR_CTRL_25                                                                          (32'h64)
`define PV_REG_PCR_CTRL_25_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_25_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_25_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_25_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_25_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_25_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_25_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_25_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_26                                                                      (32'h1001a068)
`define PV_REG_PCR_CTRL_26                                                                          (32'h68)
`define PV_REG_PCR_CTRL_26_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_26_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_26_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_26_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_26_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_26_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_26_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_26_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_27                                                                      (32'h1001a06c)
`define PV_REG_PCR_CTRL_27                                                                          (32'h6c)
`define PV_REG_PCR_CTRL_27_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_27_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_27_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_27_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_27_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_27_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_27_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_27_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_28                                                                      (32'h1001a070)
`define PV_REG_PCR_CTRL_28                                                                          (32'h70)
`define PV_REG_PCR_CTRL_28_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_28_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_28_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_28_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_28_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_28_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_28_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_28_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_29                                                                      (32'h1001a074)
`define PV_REG_PCR_CTRL_29                                                                          (32'h74)
`define PV_REG_PCR_CTRL_29_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_29_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_29_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_29_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_29_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_29_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_29_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_29_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_30                                                                      (32'h1001a078)
`define PV_REG_PCR_CTRL_30                                                                          (32'h78)
`define PV_REG_PCR_CTRL_30_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_30_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_30_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_30_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_30_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_30_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_30_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_30_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_31                                                                      (32'h1001a07c)
`define PV_REG_PCR_CTRL_31                                                                          (32'h7c)
`define PV_REG_PCR_CTRL_31_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_31_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_31_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_31_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_31_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_31_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_31_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_31_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_ENTRY_0_0                                                                    (32'h1001a600)
`define PV_REG_PCR_ENTRY_0_0                                                                        (32'h600)
`define CLP_PV_REG_PCR_ENTRY_0_1                                                                    (32'h1001a604)
`define PV_REG_PCR_ENTRY_0_1                                                                        (32'h604)
`define CLP_PV_REG_PCR_ENTRY_0_2                                                                    (32'h1001a608)
`define PV_REG_PCR_ENTRY_0_2                                                                        (32'h608)
`define CLP_PV_REG_PCR_ENTRY_0_3                                                                    (32'h1001a60c)
`define PV_REG_PCR_ENTRY_0_3                                                                        (32'h60c)
`define CLP_PV_REG_PCR_ENTRY_0_4                                                                    (32'h1001a610)
`define PV_REG_PCR_ENTRY_0_4                                                                        (32'h610)
`define CLP_PV_REG_PCR_ENTRY_0_5                                                                    (32'h1001a614)
`define PV_REG_PCR_ENTRY_0_5                                                                        (32'h614)
`define CLP_PV_REG_PCR_ENTRY_0_6                                                                    (32'h1001a618)
`define PV_REG_PCR_ENTRY_0_6                                                                        (32'h618)
`define CLP_PV_REG_PCR_ENTRY_0_7                                                                    (32'h1001a61c)
`define PV_REG_PCR_ENTRY_0_7                                                                        (32'h61c)
`define CLP_PV_REG_PCR_ENTRY_0_8                                                                    (32'h1001a620)
`define PV_REG_PCR_ENTRY_0_8                                                                        (32'h620)
`define CLP_PV_REG_PCR_ENTRY_0_9                                                                    (32'h1001a624)
`define PV_REG_PCR_ENTRY_0_9                                                                        (32'h624)
`define CLP_PV_REG_PCR_ENTRY_0_10                                                                   (32'h1001a628)
`define PV_REG_PCR_ENTRY_0_10                                                                       (32'h628)
`define CLP_PV_REG_PCR_ENTRY_0_11                                                                   (32'h1001a62c)
`define PV_REG_PCR_ENTRY_0_11                                                                       (32'h62c)
`define CLP_PV_REG_PCR_ENTRY_1_0                                                                    (32'h1001a630)
`define PV_REG_PCR_ENTRY_1_0                                                                        (32'h630)
`define CLP_PV_REG_PCR_ENTRY_1_1                                                                    (32'h1001a634)
`define PV_REG_PCR_ENTRY_1_1                                                                        (32'h634)
`define CLP_PV_REG_PCR_ENTRY_1_2                                                                    (32'h1001a638)
`define PV_REG_PCR_ENTRY_1_2                                                                        (32'h638)
`define CLP_PV_REG_PCR_ENTRY_1_3                                                                    (32'h1001a63c)
`define PV_REG_PCR_ENTRY_1_3                                                                        (32'h63c)
`define CLP_PV_REG_PCR_ENTRY_1_4                                                                    (32'h1001a640)
`define PV_REG_PCR_ENTRY_1_4                                                                        (32'h640)
`define CLP_PV_REG_PCR_ENTRY_1_5                                                                    (32'h1001a644)
`define PV_REG_PCR_ENTRY_1_5                                                                        (32'h644)
`define CLP_PV_REG_PCR_ENTRY_1_6                                                                    (32'h1001a648)
`define PV_REG_PCR_ENTRY_1_6                                                                        (32'h648)
`define CLP_PV_REG_PCR_ENTRY_1_7                                                                    (32'h1001a64c)
`define PV_REG_PCR_ENTRY_1_7                                                                        (32'h64c)
`define CLP_PV_REG_PCR_ENTRY_1_8                                                                    (32'h1001a650)
`define PV_REG_PCR_ENTRY_1_8                                                                        (32'h650)
`define CLP_PV_REG_PCR_ENTRY_1_9                                                                    (32'h1001a654)
`define PV_REG_PCR_ENTRY_1_9                                                                        (32'h654)
`define CLP_PV_REG_PCR_ENTRY_1_10                                                                   (32'h1001a658)
`define PV_REG_PCR_ENTRY_1_10                                                                       (32'h658)
`define CLP_PV_REG_PCR_ENTRY_1_11                                                                   (32'h1001a65c)
`define PV_REG_PCR_ENTRY_1_11                                                                       (32'h65c)
`define CLP_PV_REG_PCR_ENTRY_2_0                                                                    (32'h1001a660)
`define PV_REG_PCR_ENTRY_2_0                                                                        (32'h660)
`define CLP_PV_REG_PCR_ENTRY_2_1                                                                    (32'h1001a664)
`define PV_REG_PCR_ENTRY_2_1                                                                        (32'h664)
`define CLP_PV_REG_PCR_ENTRY_2_2                                                                    (32'h1001a668)
`define PV_REG_PCR_ENTRY_2_2                                                                        (32'h668)
`define CLP_PV_REG_PCR_ENTRY_2_3                                                                    (32'h1001a66c)
`define PV_REG_PCR_ENTRY_2_3                                                                        (32'h66c)
`define CLP_PV_REG_PCR_ENTRY_2_4                                                                    (32'h1001a670)
`define PV_REG_PCR_ENTRY_2_4                                                                        (32'h670)
`define CLP_PV_REG_PCR_ENTRY_2_5                                                                    (32'h1001a674)
`define PV_REG_PCR_ENTRY_2_5                                                                        (32'h674)
`define CLP_PV_REG_PCR_ENTRY_2_6                                                                    (32'h1001a678)
`define PV_REG_PCR_ENTRY_2_6                                                                        (32'h678)
`define CLP_PV_REG_PCR_ENTRY_2_7                                                                    (32'h1001a67c)
`define PV_REG_PCR_ENTRY_2_7                                                                        (32'h67c)
`define CLP_PV_REG_PCR_ENTRY_2_8                                                                    (32'h1001a680)
`define PV_REG_PCR_ENTRY_2_8                                                                        (32'h680)
`define CLP_PV_REG_PCR_ENTRY_2_9                                                                    (32'h1001a684)
`define PV_REG_PCR_ENTRY_2_9                                                                        (32'h684)
`define CLP_PV_REG_PCR_ENTRY_2_10                                                                   (32'h1001a688)
`define PV_REG_PCR_ENTRY_2_10                                                                       (32'h688)
`define CLP_PV_REG_PCR_ENTRY_2_11                                                                   (32'h1001a68c)
`define PV_REG_PCR_ENTRY_2_11                                                                       (32'h68c)
`define CLP_PV_REG_PCR_ENTRY_3_0                                                                    (32'h1001a690)
`define PV_REG_PCR_ENTRY_3_0                                                                        (32'h690)
`define CLP_PV_REG_PCR_ENTRY_3_1                                                                    (32'h1001a694)
`define PV_REG_PCR_ENTRY_3_1                                                                        (32'h694)
`define CLP_PV_REG_PCR_ENTRY_3_2                                                                    (32'h1001a698)
`define PV_REG_PCR_ENTRY_3_2                                                                        (32'h698)
`define CLP_PV_REG_PCR_ENTRY_3_3                                                                    (32'h1001a69c)
`define PV_REG_PCR_ENTRY_3_3                                                                        (32'h69c)
`define CLP_PV_REG_PCR_ENTRY_3_4                                                                    (32'h1001a6a0)
`define PV_REG_PCR_ENTRY_3_4                                                                        (32'h6a0)
`define CLP_PV_REG_PCR_ENTRY_3_5                                                                    (32'h1001a6a4)
`define PV_REG_PCR_ENTRY_3_5                                                                        (32'h6a4)
`define CLP_PV_REG_PCR_ENTRY_3_6                                                                    (32'h1001a6a8)
`define PV_REG_PCR_ENTRY_3_6                                                                        (32'h6a8)
`define CLP_PV_REG_PCR_ENTRY_3_7                                                                    (32'h1001a6ac)
`define PV_REG_PCR_ENTRY_3_7                                                                        (32'h6ac)
`define CLP_PV_REG_PCR_ENTRY_3_8                                                                    (32'h1001a6b0)
`define PV_REG_PCR_ENTRY_3_8                                                                        (32'h6b0)
`define CLP_PV_REG_PCR_ENTRY_3_9                                                                    (32'h1001a6b4)
`define PV_REG_PCR_ENTRY_3_9                                                                        (32'h6b4)
`define CLP_PV_REG_PCR_ENTRY_3_10                                                                   (32'h1001a6b8)
`define PV_REG_PCR_ENTRY_3_10                                                                       (32'h6b8)
`define CLP_PV_REG_PCR_ENTRY_3_11                                                                   (32'h1001a6bc)
`define PV_REG_PCR_ENTRY_3_11                                                                       (32'h6bc)
`define CLP_PV_REG_PCR_ENTRY_4_0                                                                    (32'h1001a6c0)
`define PV_REG_PCR_ENTRY_4_0                                                                        (32'h6c0)
`define CLP_PV_REG_PCR_ENTRY_4_1                                                                    (32'h1001a6c4)
`define PV_REG_PCR_ENTRY_4_1                                                                        (32'h6c4)
`define CLP_PV_REG_PCR_ENTRY_4_2                                                                    (32'h1001a6c8)
`define PV_REG_PCR_ENTRY_4_2                                                                        (32'h6c8)
`define CLP_PV_REG_PCR_ENTRY_4_3                                                                    (32'h1001a6cc)
`define PV_REG_PCR_ENTRY_4_3                                                                        (32'h6cc)
`define CLP_PV_REG_PCR_ENTRY_4_4                                                                    (32'h1001a6d0)
`define PV_REG_PCR_ENTRY_4_4                                                                        (32'h6d0)
`define CLP_PV_REG_PCR_ENTRY_4_5                                                                    (32'h1001a6d4)
`define PV_REG_PCR_ENTRY_4_5                                                                        (32'h6d4)
`define CLP_PV_REG_PCR_ENTRY_4_6                                                                    (32'h1001a6d8)
`define PV_REG_PCR_ENTRY_4_6                                                                        (32'h6d8)
`define CLP_PV_REG_PCR_ENTRY_4_7                                                                    (32'h1001a6dc)
`define PV_REG_PCR_ENTRY_4_7                                                                        (32'h6dc)
`define CLP_PV_REG_PCR_ENTRY_4_8                                                                    (32'h1001a6e0)
`define PV_REG_PCR_ENTRY_4_8                                                                        (32'h6e0)
`define CLP_PV_REG_PCR_ENTRY_4_9                                                                    (32'h1001a6e4)
`define PV_REG_PCR_ENTRY_4_9                                                                        (32'h6e4)
`define CLP_PV_REG_PCR_ENTRY_4_10                                                                   (32'h1001a6e8)
`define PV_REG_PCR_ENTRY_4_10                                                                       (32'h6e8)
`define CLP_PV_REG_PCR_ENTRY_4_11                                                                   (32'h1001a6ec)
`define PV_REG_PCR_ENTRY_4_11                                                                       (32'h6ec)
`define CLP_PV_REG_PCR_ENTRY_5_0                                                                    (32'h1001a6f0)
`define PV_REG_PCR_ENTRY_5_0                                                                        (32'h6f0)
`define CLP_PV_REG_PCR_ENTRY_5_1                                                                    (32'h1001a6f4)
`define PV_REG_PCR_ENTRY_5_1                                                                        (32'h6f4)
`define CLP_PV_REG_PCR_ENTRY_5_2                                                                    (32'h1001a6f8)
`define PV_REG_PCR_ENTRY_5_2                                                                        (32'h6f8)
`define CLP_PV_REG_PCR_ENTRY_5_3                                                                    (32'h1001a6fc)
`define PV_REG_PCR_ENTRY_5_3                                                                        (32'h6fc)
`define CLP_PV_REG_PCR_ENTRY_5_4                                                                    (32'h1001a700)
`define PV_REG_PCR_ENTRY_5_4                                                                        (32'h700)
`define CLP_PV_REG_PCR_ENTRY_5_5                                                                    (32'h1001a704)
`define PV_REG_PCR_ENTRY_5_5                                                                        (32'h704)
`define CLP_PV_REG_PCR_ENTRY_5_6                                                                    (32'h1001a708)
`define PV_REG_PCR_ENTRY_5_6                                                                        (32'h708)
`define CLP_PV_REG_PCR_ENTRY_5_7                                                                    (32'h1001a70c)
`define PV_REG_PCR_ENTRY_5_7                                                                        (32'h70c)
`define CLP_PV_REG_PCR_ENTRY_5_8                                                                    (32'h1001a710)
`define PV_REG_PCR_ENTRY_5_8                                                                        (32'h710)
`define CLP_PV_REG_PCR_ENTRY_5_9                                                                    (32'h1001a714)
`define PV_REG_PCR_ENTRY_5_9                                                                        (32'h714)
`define CLP_PV_REG_PCR_ENTRY_5_10                                                                   (32'h1001a718)
`define PV_REG_PCR_ENTRY_5_10                                                                       (32'h718)
`define CLP_PV_REG_PCR_ENTRY_5_11                                                                   (32'h1001a71c)
`define PV_REG_PCR_ENTRY_5_11                                                                       (32'h71c)
`define CLP_PV_REG_PCR_ENTRY_6_0                                                                    (32'h1001a720)
`define PV_REG_PCR_ENTRY_6_0                                                                        (32'h720)
`define CLP_PV_REG_PCR_ENTRY_6_1                                                                    (32'h1001a724)
`define PV_REG_PCR_ENTRY_6_1                                                                        (32'h724)
`define CLP_PV_REG_PCR_ENTRY_6_2                                                                    (32'h1001a728)
`define PV_REG_PCR_ENTRY_6_2                                                                        (32'h728)
`define CLP_PV_REG_PCR_ENTRY_6_3                                                                    (32'h1001a72c)
`define PV_REG_PCR_ENTRY_6_3                                                                        (32'h72c)
`define CLP_PV_REG_PCR_ENTRY_6_4                                                                    (32'h1001a730)
`define PV_REG_PCR_ENTRY_6_4                                                                        (32'h730)
`define CLP_PV_REG_PCR_ENTRY_6_5                                                                    (32'h1001a734)
`define PV_REG_PCR_ENTRY_6_5                                                                        (32'h734)
`define CLP_PV_REG_PCR_ENTRY_6_6                                                                    (32'h1001a738)
`define PV_REG_PCR_ENTRY_6_6                                                                        (32'h738)
`define CLP_PV_REG_PCR_ENTRY_6_7                                                                    (32'h1001a73c)
`define PV_REG_PCR_ENTRY_6_7                                                                        (32'h73c)
`define CLP_PV_REG_PCR_ENTRY_6_8                                                                    (32'h1001a740)
`define PV_REG_PCR_ENTRY_6_8                                                                        (32'h740)
`define CLP_PV_REG_PCR_ENTRY_6_9                                                                    (32'h1001a744)
`define PV_REG_PCR_ENTRY_6_9                                                                        (32'h744)
`define CLP_PV_REG_PCR_ENTRY_6_10                                                                   (32'h1001a748)
`define PV_REG_PCR_ENTRY_6_10                                                                       (32'h748)
`define CLP_PV_REG_PCR_ENTRY_6_11                                                                   (32'h1001a74c)
`define PV_REG_PCR_ENTRY_6_11                                                                       (32'h74c)
`define CLP_PV_REG_PCR_ENTRY_7_0                                                                    (32'h1001a750)
`define PV_REG_PCR_ENTRY_7_0                                                                        (32'h750)
`define CLP_PV_REG_PCR_ENTRY_7_1                                                                    (32'h1001a754)
`define PV_REG_PCR_ENTRY_7_1                                                                        (32'h754)
`define CLP_PV_REG_PCR_ENTRY_7_2                                                                    (32'h1001a758)
`define PV_REG_PCR_ENTRY_7_2                                                                        (32'h758)
`define CLP_PV_REG_PCR_ENTRY_7_3                                                                    (32'h1001a75c)
`define PV_REG_PCR_ENTRY_7_3                                                                        (32'h75c)
`define CLP_PV_REG_PCR_ENTRY_7_4                                                                    (32'h1001a760)
`define PV_REG_PCR_ENTRY_7_4                                                                        (32'h760)
`define CLP_PV_REG_PCR_ENTRY_7_5                                                                    (32'h1001a764)
`define PV_REG_PCR_ENTRY_7_5                                                                        (32'h764)
`define CLP_PV_REG_PCR_ENTRY_7_6                                                                    (32'h1001a768)
`define PV_REG_PCR_ENTRY_7_6                                                                        (32'h768)
`define CLP_PV_REG_PCR_ENTRY_7_7                                                                    (32'h1001a76c)
`define PV_REG_PCR_ENTRY_7_7                                                                        (32'h76c)
`define CLP_PV_REG_PCR_ENTRY_7_8                                                                    (32'h1001a770)
`define PV_REG_PCR_ENTRY_7_8                                                                        (32'h770)
`define CLP_PV_REG_PCR_ENTRY_7_9                                                                    (32'h1001a774)
`define PV_REG_PCR_ENTRY_7_9                                                                        (32'h774)
`define CLP_PV_REG_PCR_ENTRY_7_10                                                                   (32'h1001a778)
`define PV_REG_PCR_ENTRY_7_10                                                                       (32'h778)
`define CLP_PV_REG_PCR_ENTRY_7_11                                                                   (32'h1001a77c)
`define PV_REG_PCR_ENTRY_7_11                                                                       (32'h77c)
`define CLP_PV_REG_PCR_ENTRY_8_0                                                                    (32'h1001a780)
`define PV_REG_PCR_ENTRY_8_0                                                                        (32'h780)
`define CLP_PV_REG_PCR_ENTRY_8_1                                                                    (32'h1001a784)
`define PV_REG_PCR_ENTRY_8_1                                                                        (32'h784)
`define CLP_PV_REG_PCR_ENTRY_8_2                                                                    (32'h1001a788)
`define PV_REG_PCR_ENTRY_8_2                                                                        (32'h788)
`define CLP_PV_REG_PCR_ENTRY_8_3                                                                    (32'h1001a78c)
`define PV_REG_PCR_ENTRY_8_3                                                                        (32'h78c)
`define CLP_PV_REG_PCR_ENTRY_8_4                                                                    (32'h1001a790)
`define PV_REG_PCR_ENTRY_8_4                                                                        (32'h790)
`define CLP_PV_REG_PCR_ENTRY_8_5                                                                    (32'h1001a794)
`define PV_REG_PCR_ENTRY_8_5                                                                        (32'h794)
`define CLP_PV_REG_PCR_ENTRY_8_6                                                                    (32'h1001a798)
`define PV_REG_PCR_ENTRY_8_6                                                                        (32'h798)
`define CLP_PV_REG_PCR_ENTRY_8_7                                                                    (32'h1001a79c)
`define PV_REG_PCR_ENTRY_8_7                                                                        (32'h79c)
`define CLP_PV_REG_PCR_ENTRY_8_8                                                                    (32'h1001a7a0)
`define PV_REG_PCR_ENTRY_8_8                                                                        (32'h7a0)
`define CLP_PV_REG_PCR_ENTRY_8_9                                                                    (32'h1001a7a4)
`define PV_REG_PCR_ENTRY_8_9                                                                        (32'h7a4)
`define CLP_PV_REG_PCR_ENTRY_8_10                                                                   (32'h1001a7a8)
`define PV_REG_PCR_ENTRY_8_10                                                                       (32'h7a8)
`define CLP_PV_REG_PCR_ENTRY_8_11                                                                   (32'h1001a7ac)
`define PV_REG_PCR_ENTRY_8_11                                                                       (32'h7ac)
`define CLP_PV_REG_PCR_ENTRY_9_0                                                                    (32'h1001a7b0)
`define PV_REG_PCR_ENTRY_9_0                                                                        (32'h7b0)
`define CLP_PV_REG_PCR_ENTRY_9_1                                                                    (32'h1001a7b4)
`define PV_REG_PCR_ENTRY_9_1                                                                        (32'h7b4)
`define CLP_PV_REG_PCR_ENTRY_9_2                                                                    (32'h1001a7b8)
`define PV_REG_PCR_ENTRY_9_2                                                                        (32'h7b8)
`define CLP_PV_REG_PCR_ENTRY_9_3                                                                    (32'h1001a7bc)
`define PV_REG_PCR_ENTRY_9_3                                                                        (32'h7bc)
`define CLP_PV_REG_PCR_ENTRY_9_4                                                                    (32'h1001a7c0)
`define PV_REG_PCR_ENTRY_9_4                                                                        (32'h7c0)
`define CLP_PV_REG_PCR_ENTRY_9_5                                                                    (32'h1001a7c4)
`define PV_REG_PCR_ENTRY_9_5                                                                        (32'h7c4)
`define CLP_PV_REG_PCR_ENTRY_9_6                                                                    (32'h1001a7c8)
`define PV_REG_PCR_ENTRY_9_6                                                                        (32'h7c8)
`define CLP_PV_REG_PCR_ENTRY_9_7                                                                    (32'h1001a7cc)
`define PV_REG_PCR_ENTRY_9_7                                                                        (32'h7cc)
`define CLP_PV_REG_PCR_ENTRY_9_8                                                                    (32'h1001a7d0)
`define PV_REG_PCR_ENTRY_9_8                                                                        (32'h7d0)
`define CLP_PV_REG_PCR_ENTRY_9_9                                                                    (32'h1001a7d4)
`define PV_REG_PCR_ENTRY_9_9                                                                        (32'h7d4)
`define CLP_PV_REG_PCR_ENTRY_9_10                                                                   (32'h1001a7d8)
`define PV_REG_PCR_ENTRY_9_10                                                                       (32'h7d8)
`define CLP_PV_REG_PCR_ENTRY_9_11                                                                   (32'h1001a7dc)
`define PV_REG_PCR_ENTRY_9_11                                                                       (32'h7dc)
`define CLP_PV_REG_PCR_ENTRY_10_0                                                                   (32'h1001a7e0)
`define PV_REG_PCR_ENTRY_10_0                                                                       (32'h7e0)
`define CLP_PV_REG_PCR_ENTRY_10_1                                                                   (32'h1001a7e4)
`define PV_REG_PCR_ENTRY_10_1                                                                       (32'h7e4)
`define CLP_PV_REG_PCR_ENTRY_10_2                                                                   (32'h1001a7e8)
`define PV_REG_PCR_ENTRY_10_2                                                                       (32'h7e8)
`define CLP_PV_REG_PCR_ENTRY_10_3                                                                   (32'h1001a7ec)
`define PV_REG_PCR_ENTRY_10_3                                                                       (32'h7ec)
`define CLP_PV_REG_PCR_ENTRY_10_4                                                                   (32'h1001a7f0)
`define PV_REG_PCR_ENTRY_10_4                                                                       (32'h7f0)
`define CLP_PV_REG_PCR_ENTRY_10_5                                                                   (32'h1001a7f4)
`define PV_REG_PCR_ENTRY_10_5                                                                       (32'h7f4)
`define CLP_PV_REG_PCR_ENTRY_10_6                                                                   (32'h1001a7f8)
`define PV_REG_PCR_ENTRY_10_6                                                                       (32'h7f8)
`define CLP_PV_REG_PCR_ENTRY_10_7                                                                   (32'h1001a7fc)
`define PV_REG_PCR_ENTRY_10_7                                                                       (32'h7fc)
`define CLP_PV_REG_PCR_ENTRY_10_8                                                                   (32'h1001a800)
`define PV_REG_PCR_ENTRY_10_8                                                                       (32'h800)
`define CLP_PV_REG_PCR_ENTRY_10_9                                                                   (32'h1001a804)
`define PV_REG_PCR_ENTRY_10_9                                                                       (32'h804)
`define CLP_PV_REG_PCR_ENTRY_10_10                                                                  (32'h1001a808)
`define PV_REG_PCR_ENTRY_10_10                                                                      (32'h808)
`define CLP_PV_REG_PCR_ENTRY_10_11                                                                  (32'h1001a80c)
`define PV_REG_PCR_ENTRY_10_11                                                                      (32'h80c)
`define CLP_PV_REG_PCR_ENTRY_11_0                                                                   (32'h1001a810)
`define PV_REG_PCR_ENTRY_11_0                                                                       (32'h810)
`define CLP_PV_REG_PCR_ENTRY_11_1                                                                   (32'h1001a814)
`define PV_REG_PCR_ENTRY_11_1                                                                       (32'h814)
`define CLP_PV_REG_PCR_ENTRY_11_2                                                                   (32'h1001a818)
`define PV_REG_PCR_ENTRY_11_2                                                                       (32'h818)
`define CLP_PV_REG_PCR_ENTRY_11_3                                                                   (32'h1001a81c)
`define PV_REG_PCR_ENTRY_11_3                                                                       (32'h81c)
`define CLP_PV_REG_PCR_ENTRY_11_4                                                                   (32'h1001a820)
`define PV_REG_PCR_ENTRY_11_4                                                                       (32'h820)
`define CLP_PV_REG_PCR_ENTRY_11_5                                                                   (32'h1001a824)
`define PV_REG_PCR_ENTRY_11_5                                                                       (32'h824)
`define CLP_PV_REG_PCR_ENTRY_11_6                                                                   (32'h1001a828)
`define PV_REG_PCR_ENTRY_11_6                                                                       (32'h828)
`define CLP_PV_REG_PCR_ENTRY_11_7                                                                   (32'h1001a82c)
`define PV_REG_PCR_ENTRY_11_7                                                                       (32'h82c)
`define CLP_PV_REG_PCR_ENTRY_11_8                                                                   (32'h1001a830)
`define PV_REG_PCR_ENTRY_11_8                                                                       (32'h830)
`define CLP_PV_REG_PCR_ENTRY_11_9                                                                   (32'h1001a834)
`define PV_REG_PCR_ENTRY_11_9                                                                       (32'h834)
`define CLP_PV_REG_PCR_ENTRY_11_10                                                                  (32'h1001a838)
`define PV_REG_PCR_ENTRY_11_10                                                                      (32'h838)
`define CLP_PV_REG_PCR_ENTRY_11_11                                                                  (32'h1001a83c)
`define PV_REG_PCR_ENTRY_11_11                                                                      (32'h83c)
`define CLP_PV_REG_PCR_ENTRY_12_0                                                                   (32'h1001a840)
`define PV_REG_PCR_ENTRY_12_0                                                                       (32'h840)
`define CLP_PV_REG_PCR_ENTRY_12_1                                                                   (32'h1001a844)
`define PV_REG_PCR_ENTRY_12_1                                                                       (32'h844)
`define CLP_PV_REG_PCR_ENTRY_12_2                                                                   (32'h1001a848)
`define PV_REG_PCR_ENTRY_12_2                                                                       (32'h848)
`define CLP_PV_REG_PCR_ENTRY_12_3                                                                   (32'h1001a84c)
`define PV_REG_PCR_ENTRY_12_3                                                                       (32'h84c)
`define CLP_PV_REG_PCR_ENTRY_12_4                                                                   (32'h1001a850)
`define PV_REG_PCR_ENTRY_12_4                                                                       (32'h850)
`define CLP_PV_REG_PCR_ENTRY_12_5                                                                   (32'h1001a854)
`define PV_REG_PCR_ENTRY_12_5                                                                       (32'h854)
`define CLP_PV_REG_PCR_ENTRY_12_6                                                                   (32'h1001a858)
`define PV_REG_PCR_ENTRY_12_6                                                                       (32'h858)
`define CLP_PV_REG_PCR_ENTRY_12_7                                                                   (32'h1001a85c)
`define PV_REG_PCR_ENTRY_12_7                                                                       (32'h85c)
`define CLP_PV_REG_PCR_ENTRY_12_8                                                                   (32'h1001a860)
`define PV_REG_PCR_ENTRY_12_8                                                                       (32'h860)
`define CLP_PV_REG_PCR_ENTRY_12_9                                                                   (32'h1001a864)
`define PV_REG_PCR_ENTRY_12_9                                                                       (32'h864)
`define CLP_PV_REG_PCR_ENTRY_12_10                                                                  (32'h1001a868)
`define PV_REG_PCR_ENTRY_12_10                                                                      (32'h868)
`define CLP_PV_REG_PCR_ENTRY_12_11                                                                  (32'h1001a86c)
`define PV_REG_PCR_ENTRY_12_11                                                                      (32'h86c)
`define CLP_PV_REG_PCR_ENTRY_13_0                                                                   (32'h1001a870)
`define PV_REG_PCR_ENTRY_13_0                                                                       (32'h870)
`define CLP_PV_REG_PCR_ENTRY_13_1                                                                   (32'h1001a874)
`define PV_REG_PCR_ENTRY_13_1                                                                       (32'h874)
`define CLP_PV_REG_PCR_ENTRY_13_2                                                                   (32'h1001a878)
`define PV_REG_PCR_ENTRY_13_2                                                                       (32'h878)
`define CLP_PV_REG_PCR_ENTRY_13_3                                                                   (32'h1001a87c)
`define PV_REG_PCR_ENTRY_13_3                                                                       (32'h87c)
`define CLP_PV_REG_PCR_ENTRY_13_4                                                                   (32'h1001a880)
`define PV_REG_PCR_ENTRY_13_4                                                                       (32'h880)
`define CLP_PV_REG_PCR_ENTRY_13_5                                                                   (32'h1001a884)
`define PV_REG_PCR_ENTRY_13_5                                                                       (32'h884)
`define CLP_PV_REG_PCR_ENTRY_13_6                                                                   (32'h1001a888)
`define PV_REG_PCR_ENTRY_13_6                                                                       (32'h888)
`define CLP_PV_REG_PCR_ENTRY_13_7                                                                   (32'h1001a88c)
`define PV_REG_PCR_ENTRY_13_7                                                                       (32'h88c)
`define CLP_PV_REG_PCR_ENTRY_13_8                                                                   (32'h1001a890)
`define PV_REG_PCR_ENTRY_13_8                                                                       (32'h890)
`define CLP_PV_REG_PCR_ENTRY_13_9                                                                   (32'h1001a894)
`define PV_REG_PCR_ENTRY_13_9                                                                       (32'h894)
`define CLP_PV_REG_PCR_ENTRY_13_10                                                                  (32'h1001a898)
`define PV_REG_PCR_ENTRY_13_10                                                                      (32'h898)
`define CLP_PV_REG_PCR_ENTRY_13_11                                                                  (32'h1001a89c)
`define PV_REG_PCR_ENTRY_13_11                                                                      (32'h89c)
`define CLP_PV_REG_PCR_ENTRY_14_0                                                                   (32'h1001a8a0)
`define PV_REG_PCR_ENTRY_14_0                                                                       (32'h8a0)
`define CLP_PV_REG_PCR_ENTRY_14_1                                                                   (32'h1001a8a4)
`define PV_REG_PCR_ENTRY_14_1                                                                       (32'h8a4)
`define CLP_PV_REG_PCR_ENTRY_14_2                                                                   (32'h1001a8a8)
`define PV_REG_PCR_ENTRY_14_2                                                                       (32'h8a8)
`define CLP_PV_REG_PCR_ENTRY_14_3                                                                   (32'h1001a8ac)
`define PV_REG_PCR_ENTRY_14_3                                                                       (32'h8ac)
`define CLP_PV_REG_PCR_ENTRY_14_4                                                                   (32'h1001a8b0)
`define PV_REG_PCR_ENTRY_14_4                                                                       (32'h8b0)
`define CLP_PV_REG_PCR_ENTRY_14_5                                                                   (32'h1001a8b4)
`define PV_REG_PCR_ENTRY_14_5                                                                       (32'h8b4)
`define CLP_PV_REG_PCR_ENTRY_14_6                                                                   (32'h1001a8b8)
`define PV_REG_PCR_ENTRY_14_6                                                                       (32'h8b8)
`define CLP_PV_REG_PCR_ENTRY_14_7                                                                   (32'h1001a8bc)
`define PV_REG_PCR_ENTRY_14_7                                                                       (32'h8bc)
`define CLP_PV_REG_PCR_ENTRY_14_8                                                                   (32'h1001a8c0)
`define PV_REG_PCR_ENTRY_14_8                                                                       (32'h8c0)
`define CLP_PV_REG_PCR_ENTRY_14_9                                                                   (32'h1001a8c4)
`define PV_REG_PCR_ENTRY_14_9                                                                       (32'h8c4)
`define CLP_PV_REG_PCR_ENTRY_14_10                                                                  (32'h1001a8c8)
`define PV_REG_PCR_ENTRY_14_10                                                                      (32'h8c8)
`define CLP_PV_REG_PCR_ENTRY_14_11                                                                  (32'h1001a8cc)
`define PV_REG_PCR_ENTRY_14_11                                                                      (32'h8cc)
`define CLP_PV_REG_PCR_ENTRY_15_0                                                                   (32'h1001a8d0)
`define PV_REG_PCR_ENTRY_15_0                                                                       (32'h8d0)
`define CLP_PV_REG_PCR_ENTRY_15_1                                                                   (32'h1001a8d4)
`define PV_REG_PCR_ENTRY_15_1                                                                       (32'h8d4)
`define CLP_PV_REG_PCR_ENTRY_15_2                                                                   (32'h1001a8d8)
`define PV_REG_PCR_ENTRY_15_2                                                                       (32'h8d8)
`define CLP_PV_REG_PCR_ENTRY_15_3                                                                   (32'h1001a8dc)
`define PV_REG_PCR_ENTRY_15_3                                                                       (32'h8dc)
`define CLP_PV_REG_PCR_ENTRY_15_4                                                                   (32'h1001a8e0)
`define PV_REG_PCR_ENTRY_15_4                                                                       (32'h8e0)
`define CLP_PV_REG_PCR_ENTRY_15_5                                                                   (32'h1001a8e4)
`define PV_REG_PCR_ENTRY_15_5                                                                       (32'h8e4)
`define CLP_PV_REG_PCR_ENTRY_15_6                                                                   (32'h1001a8e8)
`define PV_REG_PCR_ENTRY_15_6                                                                       (32'h8e8)
`define CLP_PV_REG_PCR_ENTRY_15_7                                                                   (32'h1001a8ec)
`define PV_REG_PCR_ENTRY_15_7                                                                       (32'h8ec)
`define CLP_PV_REG_PCR_ENTRY_15_8                                                                   (32'h1001a8f0)
`define PV_REG_PCR_ENTRY_15_8                                                                       (32'h8f0)
`define CLP_PV_REG_PCR_ENTRY_15_9                                                                   (32'h1001a8f4)
`define PV_REG_PCR_ENTRY_15_9                                                                       (32'h8f4)
`define CLP_PV_REG_PCR_ENTRY_15_10                                                                  (32'h1001a8f8)
`define PV_REG_PCR_ENTRY_15_10                                                                      (32'h8f8)
`define CLP_PV_REG_PCR_ENTRY_15_11                                                                  (32'h1001a8fc)
`define PV_REG_PCR_ENTRY_15_11                                                                      (32'h8fc)
`define CLP_PV_REG_PCR_ENTRY_16_0                                                                   (32'h1001a900)
`define PV_REG_PCR_ENTRY_16_0                                                                       (32'h900)
`define CLP_PV_REG_PCR_ENTRY_16_1                                                                   (32'h1001a904)
`define PV_REG_PCR_ENTRY_16_1                                                                       (32'h904)
`define CLP_PV_REG_PCR_ENTRY_16_2                                                                   (32'h1001a908)
`define PV_REG_PCR_ENTRY_16_2                                                                       (32'h908)
`define CLP_PV_REG_PCR_ENTRY_16_3                                                                   (32'h1001a90c)
`define PV_REG_PCR_ENTRY_16_3                                                                       (32'h90c)
`define CLP_PV_REG_PCR_ENTRY_16_4                                                                   (32'h1001a910)
`define PV_REG_PCR_ENTRY_16_4                                                                       (32'h910)
`define CLP_PV_REG_PCR_ENTRY_16_5                                                                   (32'h1001a914)
`define PV_REG_PCR_ENTRY_16_5                                                                       (32'h914)
`define CLP_PV_REG_PCR_ENTRY_16_6                                                                   (32'h1001a918)
`define PV_REG_PCR_ENTRY_16_6                                                                       (32'h918)
`define CLP_PV_REG_PCR_ENTRY_16_7                                                                   (32'h1001a91c)
`define PV_REG_PCR_ENTRY_16_7                                                                       (32'h91c)
`define CLP_PV_REG_PCR_ENTRY_16_8                                                                   (32'h1001a920)
`define PV_REG_PCR_ENTRY_16_8                                                                       (32'h920)
`define CLP_PV_REG_PCR_ENTRY_16_9                                                                   (32'h1001a924)
`define PV_REG_PCR_ENTRY_16_9                                                                       (32'h924)
`define CLP_PV_REG_PCR_ENTRY_16_10                                                                  (32'h1001a928)
`define PV_REG_PCR_ENTRY_16_10                                                                      (32'h928)
`define CLP_PV_REG_PCR_ENTRY_16_11                                                                  (32'h1001a92c)
`define PV_REG_PCR_ENTRY_16_11                                                                      (32'h92c)
`define CLP_PV_REG_PCR_ENTRY_17_0                                                                   (32'h1001a930)
`define PV_REG_PCR_ENTRY_17_0                                                                       (32'h930)
`define CLP_PV_REG_PCR_ENTRY_17_1                                                                   (32'h1001a934)
`define PV_REG_PCR_ENTRY_17_1                                                                       (32'h934)
`define CLP_PV_REG_PCR_ENTRY_17_2                                                                   (32'h1001a938)
`define PV_REG_PCR_ENTRY_17_2                                                                       (32'h938)
`define CLP_PV_REG_PCR_ENTRY_17_3                                                                   (32'h1001a93c)
`define PV_REG_PCR_ENTRY_17_3                                                                       (32'h93c)
`define CLP_PV_REG_PCR_ENTRY_17_4                                                                   (32'h1001a940)
`define PV_REG_PCR_ENTRY_17_4                                                                       (32'h940)
`define CLP_PV_REG_PCR_ENTRY_17_5                                                                   (32'h1001a944)
`define PV_REG_PCR_ENTRY_17_5                                                                       (32'h944)
`define CLP_PV_REG_PCR_ENTRY_17_6                                                                   (32'h1001a948)
`define PV_REG_PCR_ENTRY_17_6                                                                       (32'h948)
`define CLP_PV_REG_PCR_ENTRY_17_7                                                                   (32'h1001a94c)
`define PV_REG_PCR_ENTRY_17_7                                                                       (32'h94c)
`define CLP_PV_REG_PCR_ENTRY_17_8                                                                   (32'h1001a950)
`define PV_REG_PCR_ENTRY_17_8                                                                       (32'h950)
`define CLP_PV_REG_PCR_ENTRY_17_9                                                                   (32'h1001a954)
`define PV_REG_PCR_ENTRY_17_9                                                                       (32'h954)
`define CLP_PV_REG_PCR_ENTRY_17_10                                                                  (32'h1001a958)
`define PV_REG_PCR_ENTRY_17_10                                                                      (32'h958)
`define CLP_PV_REG_PCR_ENTRY_17_11                                                                  (32'h1001a95c)
`define PV_REG_PCR_ENTRY_17_11                                                                      (32'h95c)
`define CLP_PV_REG_PCR_ENTRY_18_0                                                                   (32'h1001a960)
`define PV_REG_PCR_ENTRY_18_0                                                                       (32'h960)
`define CLP_PV_REG_PCR_ENTRY_18_1                                                                   (32'h1001a964)
`define PV_REG_PCR_ENTRY_18_1                                                                       (32'h964)
`define CLP_PV_REG_PCR_ENTRY_18_2                                                                   (32'h1001a968)
`define PV_REG_PCR_ENTRY_18_2                                                                       (32'h968)
`define CLP_PV_REG_PCR_ENTRY_18_3                                                                   (32'h1001a96c)
`define PV_REG_PCR_ENTRY_18_3                                                                       (32'h96c)
`define CLP_PV_REG_PCR_ENTRY_18_4                                                                   (32'h1001a970)
`define PV_REG_PCR_ENTRY_18_4                                                                       (32'h970)
`define CLP_PV_REG_PCR_ENTRY_18_5                                                                   (32'h1001a974)
`define PV_REG_PCR_ENTRY_18_5                                                                       (32'h974)
`define CLP_PV_REG_PCR_ENTRY_18_6                                                                   (32'h1001a978)
`define PV_REG_PCR_ENTRY_18_6                                                                       (32'h978)
`define CLP_PV_REG_PCR_ENTRY_18_7                                                                   (32'h1001a97c)
`define PV_REG_PCR_ENTRY_18_7                                                                       (32'h97c)
`define CLP_PV_REG_PCR_ENTRY_18_8                                                                   (32'h1001a980)
`define PV_REG_PCR_ENTRY_18_8                                                                       (32'h980)
`define CLP_PV_REG_PCR_ENTRY_18_9                                                                   (32'h1001a984)
`define PV_REG_PCR_ENTRY_18_9                                                                       (32'h984)
`define CLP_PV_REG_PCR_ENTRY_18_10                                                                  (32'h1001a988)
`define PV_REG_PCR_ENTRY_18_10                                                                      (32'h988)
`define CLP_PV_REG_PCR_ENTRY_18_11                                                                  (32'h1001a98c)
`define PV_REG_PCR_ENTRY_18_11                                                                      (32'h98c)
`define CLP_PV_REG_PCR_ENTRY_19_0                                                                   (32'h1001a990)
`define PV_REG_PCR_ENTRY_19_0                                                                       (32'h990)
`define CLP_PV_REG_PCR_ENTRY_19_1                                                                   (32'h1001a994)
`define PV_REG_PCR_ENTRY_19_1                                                                       (32'h994)
`define CLP_PV_REG_PCR_ENTRY_19_2                                                                   (32'h1001a998)
`define PV_REG_PCR_ENTRY_19_2                                                                       (32'h998)
`define CLP_PV_REG_PCR_ENTRY_19_3                                                                   (32'h1001a99c)
`define PV_REG_PCR_ENTRY_19_3                                                                       (32'h99c)
`define CLP_PV_REG_PCR_ENTRY_19_4                                                                   (32'h1001a9a0)
`define PV_REG_PCR_ENTRY_19_4                                                                       (32'h9a0)
`define CLP_PV_REG_PCR_ENTRY_19_5                                                                   (32'h1001a9a4)
`define PV_REG_PCR_ENTRY_19_5                                                                       (32'h9a4)
`define CLP_PV_REG_PCR_ENTRY_19_6                                                                   (32'h1001a9a8)
`define PV_REG_PCR_ENTRY_19_6                                                                       (32'h9a8)
`define CLP_PV_REG_PCR_ENTRY_19_7                                                                   (32'h1001a9ac)
`define PV_REG_PCR_ENTRY_19_7                                                                       (32'h9ac)
`define CLP_PV_REG_PCR_ENTRY_19_8                                                                   (32'h1001a9b0)
`define PV_REG_PCR_ENTRY_19_8                                                                       (32'h9b0)
`define CLP_PV_REG_PCR_ENTRY_19_9                                                                   (32'h1001a9b4)
`define PV_REG_PCR_ENTRY_19_9                                                                       (32'h9b4)
`define CLP_PV_REG_PCR_ENTRY_19_10                                                                  (32'h1001a9b8)
`define PV_REG_PCR_ENTRY_19_10                                                                      (32'h9b8)
`define CLP_PV_REG_PCR_ENTRY_19_11                                                                  (32'h1001a9bc)
`define PV_REG_PCR_ENTRY_19_11                                                                      (32'h9bc)
`define CLP_PV_REG_PCR_ENTRY_20_0                                                                   (32'h1001a9c0)
`define PV_REG_PCR_ENTRY_20_0                                                                       (32'h9c0)
`define CLP_PV_REG_PCR_ENTRY_20_1                                                                   (32'h1001a9c4)
`define PV_REG_PCR_ENTRY_20_1                                                                       (32'h9c4)
`define CLP_PV_REG_PCR_ENTRY_20_2                                                                   (32'h1001a9c8)
`define PV_REG_PCR_ENTRY_20_2                                                                       (32'h9c8)
`define CLP_PV_REG_PCR_ENTRY_20_3                                                                   (32'h1001a9cc)
`define PV_REG_PCR_ENTRY_20_3                                                                       (32'h9cc)
`define CLP_PV_REG_PCR_ENTRY_20_4                                                                   (32'h1001a9d0)
`define PV_REG_PCR_ENTRY_20_4                                                                       (32'h9d0)
`define CLP_PV_REG_PCR_ENTRY_20_5                                                                   (32'h1001a9d4)
`define PV_REG_PCR_ENTRY_20_5                                                                       (32'h9d4)
`define CLP_PV_REG_PCR_ENTRY_20_6                                                                   (32'h1001a9d8)
`define PV_REG_PCR_ENTRY_20_6                                                                       (32'h9d8)
`define CLP_PV_REG_PCR_ENTRY_20_7                                                                   (32'h1001a9dc)
`define PV_REG_PCR_ENTRY_20_7                                                                       (32'h9dc)
`define CLP_PV_REG_PCR_ENTRY_20_8                                                                   (32'h1001a9e0)
`define PV_REG_PCR_ENTRY_20_8                                                                       (32'h9e0)
`define CLP_PV_REG_PCR_ENTRY_20_9                                                                   (32'h1001a9e4)
`define PV_REG_PCR_ENTRY_20_9                                                                       (32'h9e4)
`define CLP_PV_REG_PCR_ENTRY_20_10                                                                  (32'h1001a9e8)
`define PV_REG_PCR_ENTRY_20_10                                                                      (32'h9e8)
`define CLP_PV_REG_PCR_ENTRY_20_11                                                                  (32'h1001a9ec)
`define PV_REG_PCR_ENTRY_20_11                                                                      (32'h9ec)
`define CLP_PV_REG_PCR_ENTRY_21_0                                                                   (32'h1001a9f0)
`define PV_REG_PCR_ENTRY_21_0                                                                       (32'h9f0)
`define CLP_PV_REG_PCR_ENTRY_21_1                                                                   (32'h1001a9f4)
`define PV_REG_PCR_ENTRY_21_1                                                                       (32'h9f4)
`define CLP_PV_REG_PCR_ENTRY_21_2                                                                   (32'h1001a9f8)
`define PV_REG_PCR_ENTRY_21_2                                                                       (32'h9f8)
`define CLP_PV_REG_PCR_ENTRY_21_3                                                                   (32'h1001a9fc)
`define PV_REG_PCR_ENTRY_21_3                                                                       (32'h9fc)
`define CLP_PV_REG_PCR_ENTRY_21_4                                                                   (32'h1001aa00)
`define PV_REG_PCR_ENTRY_21_4                                                                       (32'ha00)
`define CLP_PV_REG_PCR_ENTRY_21_5                                                                   (32'h1001aa04)
`define PV_REG_PCR_ENTRY_21_5                                                                       (32'ha04)
`define CLP_PV_REG_PCR_ENTRY_21_6                                                                   (32'h1001aa08)
`define PV_REG_PCR_ENTRY_21_6                                                                       (32'ha08)
`define CLP_PV_REG_PCR_ENTRY_21_7                                                                   (32'h1001aa0c)
`define PV_REG_PCR_ENTRY_21_7                                                                       (32'ha0c)
`define CLP_PV_REG_PCR_ENTRY_21_8                                                                   (32'h1001aa10)
`define PV_REG_PCR_ENTRY_21_8                                                                       (32'ha10)
`define CLP_PV_REG_PCR_ENTRY_21_9                                                                   (32'h1001aa14)
`define PV_REG_PCR_ENTRY_21_9                                                                       (32'ha14)
`define CLP_PV_REG_PCR_ENTRY_21_10                                                                  (32'h1001aa18)
`define PV_REG_PCR_ENTRY_21_10                                                                      (32'ha18)
`define CLP_PV_REG_PCR_ENTRY_21_11                                                                  (32'h1001aa1c)
`define PV_REG_PCR_ENTRY_21_11                                                                      (32'ha1c)
`define CLP_PV_REG_PCR_ENTRY_22_0                                                                   (32'h1001aa20)
`define PV_REG_PCR_ENTRY_22_0                                                                       (32'ha20)
`define CLP_PV_REG_PCR_ENTRY_22_1                                                                   (32'h1001aa24)
`define PV_REG_PCR_ENTRY_22_1                                                                       (32'ha24)
`define CLP_PV_REG_PCR_ENTRY_22_2                                                                   (32'h1001aa28)
`define PV_REG_PCR_ENTRY_22_2                                                                       (32'ha28)
`define CLP_PV_REG_PCR_ENTRY_22_3                                                                   (32'h1001aa2c)
`define PV_REG_PCR_ENTRY_22_3                                                                       (32'ha2c)
`define CLP_PV_REG_PCR_ENTRY_22_4                                                                   (32'h1001aa30)
`define PV_REG_PCR_ENTRY_22_4                                                                       (32'ha30)
`define CLP_PV_REG_PCR_ENTRY_22_5                                                                   (32'h1001aa34)
`define PV_REG_PCR_ENTRY_22_5                                                                       (32'ha34)
`define CLP_PV_REG_PCR_ENTRY_22_6                                                                   (32'h1001aa38)
`define PV_REG_PCR_ENTRY_22_6                                                                       (32'ha38)
`define CLP_PV_REG_PCR_ENTRY_22_7                                                                   (32'h1001aa3c)
`define PV_REG_PCR_ENTRY_22_7                                                                       (32'ha3c)
`define CLP_PV_REG_PCR_ENTRY_22_8                                                                   (32'h1001aa40)
`define PV_REG_PCR_ENTRY_22_8                                                                       (32'ha40)
`define CLP_PV_REG_PCR_ENTRY_22_9                                                                   (32'h1001aa44)
`define PV_REG_PCR_ENTRY_22_9                                                                       (32'ha44)
`define CLP_PV_REG_PCR_ENTRY_22_10                                                                  (32'h1001aa48)
`define PV_REG_PCR_ENTRY_22_10                                                                      (32'ha48)
`define CLP_PV_REG_PCR_ENTRY_22_11                                                                  (32'h1001aa4c)
`define PV_REG_PCR_ENTRY_22_11                                                                      (32'ha4c)
`define CLP_PV_REG_PCR_ENTRY_23_0                                                                   (32'h1001aa50)
`define PV_REG_PCR_ENTRY_23_0                                                                       (32'ha50)
`define CLP_PV_REG_PCR_ENTRY_23_1                                                                   (32'h1001aa54)
`define PV_REG_PCR_ENTRY_23_1                                                                       (32'ha54)
`define CLP_PV_REG_PCR_ENTRY_23_2                                                                   (32'h1001aa58)
`define PV_REG_PCR_ENTRY_23_2                                                                       (32'ha58)
`define CLP_PV_REG_PCR_ENTRY_23_3                                                                   (32'h1001aa5c)
`define PV_REG_PCR_ENTRY_23_3                                                                       (32'ha5c)
`define CLP_PV_REG_PCR_ENTRY_23_4                                                                   (32'h1001aa60)
`define PV_REG_PCR_ENTRY_23_4                                                                       (32'ha60)
`define CLP_PV_REG_PCR_ENTRY_23_5                                                                   (32'h1001aa64)
`define PV_REG_PCR_ENTRY_23_5                                                                       (32'ha64)
`define CLP_PV_REG_PCR_ENTRY_23_6                                                                   (32'h1001aa68)
`define PV_REG_PCR_ENTRY_23_6                                                                       (32'ha68)
`define CLP_PV_REG_PCR_ENTRY_23_7                                                                   (32'h1001aa6c)
`define PV_REG_PCR_ENTRY_23_7                                                                       (32'ha6c)
`define CLP_PV_REG_PCR_ENTRY_23_8                                                                   (32'h1001aa70)
`define PV_REG_PCR_ENTRY_23_8                                                                       (32'ha70)
`define CLP_PV_REG_PCR_ENTRY_23_9                                                                   (32'h1001aa74)
`define PV_REG_PCR_ENTRY_23_9                                                                       (32'ha74)
`define CLP_PV_REG_PCR_ENTRY_23_10                                                                  (32'h1001aa78)
`define PV_REG_PCR_ENTRY_23_10                                                                      (32'ha78)
`define CLP_PV_REG_PCR_ENTRY_23_11                                                                  (32'h1001aa7c)
`define PV_REG_PCR_ENTRY_23_11                                                                      (32'ha7c)
`define CLP_PV_REG_PCR_ENTRY_24_0                                                                   (32'h1001aa80)
`define PV_REG_PCR_ENTRY_24_0                                                                       (32'ha80)
`define CLP_PV_REG_PCR_ENTRY_24_1                                                                   (32'h1001aa84)
`define PV_REG_PCR_ENTRY_24_1                                                                       (32'ha84)
`define CLP_PV_REG_PCR_ENTRY_24_2                                                                   (32'h1001aa88)
`define PV_REG_PCR_ENTRY_24_2                                                                       (32'ha88)
`define CLP_PV_REG_PCR_ENTRY_24_3                                                                   (32'h1001aa8c)
`define PV_REG_PCR_ENTRY_24_3                                                                       (32'ha8c)
`define CLP_PV_REG_PCR_ENTRY_24_4                                                                   (32'h1001aa90)
`define PV_REG_PCR_ENTRY_24_4                                                                       (32'ha90)
`define CLP_PV_REG_PCR_ENTRY_24_5                                                                   (32'h1001aa94)
`define PV_REG_PCR_ENTRY_24_5                                                                       (32'ha94)
`define CLP_PV_REG_PCR_ENTRY_24_6                                                                   (32'h1001aa98)
`define PV_REG_PCR_ENTRY_24_6                                                                       (32'ha98)
`define CLP_PV_REG_PCR_ENTRY_24_7                                                                   (32'h1001aa9c)
`define PV_REG_PCR_ENTRY_24_7                                                                       (32'ha9c)
`define CLP_PV_REG_PCR_ENTRY_24_8                                                                   (32'h1001aaa0)
`define PV_REG_PCR_ENTRY_24_8                                                                       (32'haa0)
`define CLP_PV_REG_PCR_ENTRY_24_9                                                                   (32'h1001aaa4)
`define PV_REG_PCR_ENTRY_24_9                                                                       (32'haa4)
`define CLP_PV_REG_PCR_ENTRY_24_10                                                                  (32'h1001aaa8)
`define PV_REG_PCR_ENTRY_24_10                                                                      (32'haa8)
`define CLP_PV_REG_PCR_ENTRY_24_11                                                                  (32'h1001aaac)
`define PV_REG_PCR_ENTRY_24_11                                                                      (32'haac)
`define CLP_PV_REG_PCR_ENTRY_25_0                                                                   (32'h1001aab0)
`define PV_REG_PCR_ENTRY_25_0                                                                       (32'hab0)
`define CLP_PV_REG_PCR_ENTRY_25_1                                                                   (32'h1001aab4)
`define PV_REG_PCR_ENTRY_25_1                                                                       (32'hab4)
`define CLP_PV_REG_PCR_ENTRY_25_2                                                                   (32'h1001aab8)
`define PV_REG_PCR_ENTRY_25_2                                                                       (32'hab8)
`define CLP_PV_REG_PCR_ENTRY_25_3                                                                   (32'h1001aabc)
`define PV_REG_PCR_ENTRY_25_3                                                                       (32'habc)
`define CLP_PV_REG_PCR_ENTRY_25_4                                                                   (32'h1001aac0)
`define PV_REG_PCR_ENTRY_25_4                                                                       (32'hac0)
`define CLP_PV_REG_PCR_ENTRY_25_5                                                                   (32'h1001aac4)
`define PV_REG_PCR_ENTRY_25_5                                                                       (32'hac4)
`define CLP_PV_REG_PCR_ENTRY_25_6                                                                   (32'h1001aac8)
`define PV_REG_PCR_ENTRY_25_6                                                                       (32'hac8)
`define CLP_PV_REG_PCR_ENTRY_25_7                                                                   (32'h1001aacc)
`define PV_REG_PCR_ENTRY_25_7                                                                       (32'hacc)
`define CLP_PV_REG_PCR_ENTRY_25_8                                                                   (32'h1001aad0)
`define PV_REG_PCR_ENTRY_25_8                                                                       (32'had0)
`define CLP_PV_REG_PCR_ENTRY_25_9                                                                   (32'h1001aad4)
`define PV_REG_PCR_ENTRY_25_9                                                                       (32'had4)
`define CLP_PV_REG_PCR_ENTRY_25_10                                                                  (32'h1001aad8)
`define PV_REG_PCR_ENTRY_25_10                                                                      (32'had8)
`define CLP_PV_REG_PCR_ENTRY_25_11                                                                  (32'h1001aadc)
`define PV_REG_PCR_ENTRY_25_11                                                                      (32'hadc)
`define CLP_PV_REG_PCR_ENTRY_26_0                                                                   (32'h1001aae0)
`define PV_REG_PCR_ENTRY_26_0                                                                       (32'hae0)
`define CLP_PV_REG_PCR_ENTRY_26_1                                                                   (32'h1001aae4)
`define PV_REG_PCR_ENTRY_26_1                                                                       (32'hae4)
`define CLP_PV_REG_PCR_ENTRY_26_2                                                                   (32'h1001aae8)
`define PV_REG_PCR_ENTRY_26_2                                                                       (32'hae8)
`define CLP_PV_REG_PCR_ENTRY_26_3                                                                   (32'h1001aaec)
`define PV_REG_PCR_ENTRY_26_3                                                                       (32'haec)
`define CLP_PV_REG_PCR_ENTRY_26_4                                                                   (32'h1001aaf0)
`define PV_REG_PCR_ENTRY_26_4                                                                       (32'haf0)
`define CLP_PV_REG_PCR_ENTRY_26_5                                                                   (32'h1001aaf4)
`define PV_REG_PCR_ENTRY_26_5                                                                       (32'haf4)
`define CLP_PV_REG_PCR_ENTRY_26_6                                                                   (32'h1001aaf8)
`define PV_REG_PCR_ENTRY_26_6                                                                       (32'haf8)
`define CLP_PV_REG_PCR_ENTRY_26_7                                                                   (32'h1001aafc)
`define PV_REG_PCR_ENTRY_26_7                                                                       (32'hafc)
`define CLP_PV_REG_PCR_ENTRY_26_8                                                                   (32'h1001ab00)
`define PV_REG_PCR_ENTRY_26_8                                                                       (32'hb00)
`define CLP_PV_REG_PCR_ENTRY_26_9                                                                   (32'h1001ab04)
`define PV_REG_PCR_ENTRY_26_9                                                                       (32'hb04)
`define CLP_PV_REG_PCR_ENTRY_26_10                                                                  (32'h1001ab08)
`define PV_REG_PCR_ENTRY_26_10                                                                      (32'hb08)
`define CLP_PV_REG_PCR_ENTRY_26_11                                                                  (32'h1001ab0c)
`define PV_REG_PCR_ENTRY_26_11                                                                      (32'hb0c)
`define CLP_PV_REG_PCR_ENTRY_27_0                                                                   (32'h1001ab10)
`define PV_REG_PCR_ENTRY_27_0                                                                       (32'hb10)
`define CLP_PV_REG_PCR_ENTRY_27_1                                                                   (32'h1001ab14)
`define PV_REG_PCR_ENTRY_27_1                                                                       (32'hb14)
`define CLP_PV_REG_PCR_ENTRY_27_2                                                                   (32'h1001ab18)
`define PV_REG_PCR_ENTRY_27_2                                                                       (32'hb18)
`define CLP_PV_REG_PCR_ENTRY_27_3                                                                   (32'h1001ab1c)
`define PV_REG_PCR_ENTRY_27_3                                                                       (32'hb1c)
`define CLP_PV_REG_PCR_ENTRY_27_4                                                                   (32'h1001ab20)
`define PV_REG_PCR_ENTRY_27_4                                                                       (32'hb20)
`define CLP_PV_REG_PCR_ENTRY_27_5                                                                   (32'h1001ab24)
`define PV_REG_PCR_ENTRY_27_5                                                                       (32'hb24)
`define CLP_PV_REG_PCR_ENTRY_27_6                                                                   (32'h1001ab28)
`define PV_REG_PCR_ENTRY_27_6                                                                       (32'hb28)
`define CLP_PV_REG_PCR_ENTRY_27_7                                                                   (32'h1001ab2c)
`define PV_REG_PCR_ENTRY_27_7                                                                       (32'hb2c)
`define CLP_PV_REG_PCR_ENTRY_27_8                                                                   (32'h1001ab30)
`define PV_REG_PCR_ENTRY_27_8                                                                       (32'hb30)
`define CLP_PV_REG_PCR_ENTRY_27_9                                                                   (32'h1001ab34)
`define PV_REG_PCR_ENTRY_27_9                                                                       (32'hb34)
`define CLP_PV_REG_PCR_ENTRY_27_10                                                                  (32'h1001ab38)
`define PV_REG_PCR_ENTRY_27_10                                                                      (32'hb38)
`define CLP_PV_REG_PCR_ENTRY_27_11                                                                  (32'h1001ab3c)
`define PV_REG_PCR_ENTRY_27_11                                                                      (32'hb3c)
`define CLP_PV_REG_PCR_ENTRY_28_0                                                                   (32'h1001ab40)
`define PV_REG_PCR_ENTRY_28_0                                                                       (32'hb40)
`define CLP_PV_REG_PCR_ENTRY_28_1                                                                   (32'h1001ab44)
`define PV_REG_PCR_ENTRY_28_1                                                                       (32'hb44)
`define CLP_PV_REG_PCR_ENTRY_28_2                                                                   (32'h1001ab48)
`define PV_REG_PCR_ENTRY_28_2                                                                       (32'hb48)
`define CLP_PV_REG_PCR_ENTRY_28_3                                                                   (32'h1001ab4c)
`define PV_REG_PCR_ENTRY_28_3                                                                       (32'hb4c)
`define CLP_PV_REG_PCR_ENTRY_28_4                                                                   (32'h1001ab50)
`define PV_REG_PCR_ENTRY_28_4                                                                       (32'hb50)
`define CLP_PV_REG_PCR_ENTRY_28_5                                                                   (32'h1001ab54)
`define PV_REG_PCR_ENTRY_28_5                                                                       (32'hb54)
`define CLP_PV_REG_PCR_ENTRY_28_6                                                                   (32'h1001ab58)
`define PV_REG_PCR_ENTRY_28_6                                                                       (32'hb58)
`define CLP_PV_REG_PCR_ENTRY_28_7                                                                   (32'h1001ab5c)
`define PV_REG_PCR_ENTRY_28_7                                                                       (32'hb5c)
`define CLP_PV_REG_PCR_ENTRY_28_8                                                                   (32'h1001ab60)
`define PV_REG_PCR_ENTRY_28_8                                                                       (32'hb60)
`define CLP_PV_REG_PCR_ENTRY_28_9                                                                   (32'h1001ab64)
`define PV_REG_PCR_ENTRY_28_9                                                                       (32'hb64)
`define CLP_PV_REG_PCR_ENTRY_28_10                                                                  (32'h1001ab68)
`define PV_REG_PCR_ENTRY_28_10                                                                      (32'hb68)
`define CLP_PV_REG_PCR_ENTRY_28_11                                                                  (32'h1001ab6c)
`define PV_REG_PCR_ENTRY_28_11                                                                      (32'hb6c)
`define CLP_PV_REG_PCR_ENTRY_29_0                                                                   (32'h1001ab70)
`define PV_REG_PCR_ENTRY_29_0                                                                       (32'hb70)
`define CLP_PV_REG_PCR_ENTRY_29_1                                                                   (32'h1001ab74)
`define PV_REG_PCR_ENTRY_29_1                                                                       (32'hb74)
`define CLP_PV_REG_PCR_ENTRY_29_2                                                                   (32'h1001ab78)
`define PV_REG_PCR_ENTRY_29_2                                                                       (32'hb78)
`define CLP_PV_REG_PCR_ENTRY_29_3                                                                   (32'h1001ab7c)
`define PV_REG_PCR_ENTRY_29_3                                                                       (32'hb7c)
`define CLP_PV_REG_PCR_ENTRY_29_4                                                                   (32'h1001ab80)
`define PV_REG_PCR_ENTRY_29_4                                                                       (32'hb80)
`define CLP_PV_REG_PCR_ENTRY_29_5                                                                   (32'h1001ab84)
`define PV_REG_PCR_ENTRY_29_5                                                                       (32'hb84)
`define CLP_PV_REG_PCR_ENTRY_29_6                                                                   (32'h1001ab88)
`define PV_REG_PCR_ENTRY_29_6                                                                       (32'hb88)
`define CLP_PV_REG_PCR_ENTRY_29_7                                                                   (32'h1001ab8c)
`define PV_REG_PCR_ENTRY_29_7                                                                       (32'hb8c)
`define CLP_PV_REG_PCR_ENTRY_29_8                                                                   (32'h1001ab90)
`define PV_REG_PCR_ENTRY_29_8                                                                       (32'hb90)
`define CLP_PV_REG_PCR_ENTRY_29_9                                                                   (32'h1001ab94)
`define PV_REG_PCR_ENTRY_29_9                                                                       (32'hb94)
`define CLP_PV_REG_PCR_ENTRY_29_10                                                                  (32'h1001ab98)
`define PV_REG_PCR_ENTRY_29_10                                                                      (32'hb98)
`define CLP_PV_REG_PCR_ENTRY_29_11                                                                  (32'h1001ab9c)
`define PV_REG_PCR_ENTRY_29_11                                                                      (32'hb9c)
`define CLP_PV_REG_PCR_ENTRY_30_0                                                                   (32'h1001aba0)
`define PV_REG_PCR_ENTRY_30_0                                                                       (32'hba0)
`define CLP_PV_REG_PCR_ENTRY_30_1                                                                   (32'h1001aba4)
`define PV_REG_PCR_ENTRY_30_1                                                                       (32'hba4)
`define CLP_PV_REG_PCR_ENTRY_30_2                                                                   (32'h1001aba8)
`define PV_REG_PCR_ENTRY_30_2                                                                       (32'hba8)
`define CLP_PV_REG_PCR_ENTRY_30_3                                                                   (32'h1001abac)
`define PV_REG_PCR_ENTRY_30_3                                                                       (32'hbac)
`define CLP_PV_REG_PCR_ENTRY_30_4                                                                   (32'h1001abb0)
`define PV_REG_PCR_ENTRY_30_4                                                                       (32'hbb0)
`define CLP_PV_REG_PCR_ENTRY_30_5                                                                   (32'h1001abb4)
`define PV_REG_PCR_ENTRY_30_5                                                                       (32'hbb4)
`define CLP_PV_REG_PCR_ENTRY_30_6                                                                   (32'h1001abb8)
`define PV_REG_PCR_ENTRY_30_6                                                                       (32'hbb8)
`define CLP_PV_REG_PCR_ENTRY_30_7                                                                   (32'h1001abbc)
`define PV_REG_PCR_ENTRY_30_7                                                                       (32'hbbc)
`define CLP_PV_REG_PCR_ENTRY_30_8                                                                   (32'h1001abc0)
`define PV_REG_PCR_ENTRY_30_8                                                                       (32'hbc0)
`define CLP_PV_REG_PCR_ENTRY_30_9                                                                   (32'h1001abc4)
`define PV_REG_PCR_ENTRY_30_9                                                                       (32'hbc4)
`define CLP_PV_REG_PCR_ENTRY_30_10                                                                  (32'h1001abc8)
`define PV_REG_PCR_ENTRY_30_10                                                                      (32'hbc8)
`define CLP_PV_REG_PCR_ENTRY_30_11                                                                  (32'h1001abcc)
`define PV_REG_PCR_ENTRY_30_11                                                                      (32'hbcc)
`define CLP_PV_REG_PCR_ENTRY_31_0                                                                   (32'h1001abd0)
`define PV_REG_PCR_ENTRY_31_0                                                                       (32'hbd0)
`define CLP_PV_REG_PCR_ENTRY_31_1                                                                   (32'h1001abd4)
`define PV_REG_PCR_ENTRY_31_1                                                                       (32'hbd4)
`define CLP_PV_REG_PCR_ENTRY_31_2                                                                   (32'h1001abd8)
`define PV_REG_PCR_ENTRY_31_2                                                                       (32'hbd8)
`define CLP_PV_REG_PCR_ENTRY_31_3                                                                   (32'h1001abdc)
`define PV_REG_PCR_ENTRY_31_3                                                                       (32'hbdc)
`define CLP_PV_REG_PCR_ENTRY_31_4                                                                   (32'h1001abe0)
`define PV_REG_PCR_ENTRY_31_4                                                                       (32'hbe0)
`define CLP_PV_REG_PCR_ENTRY_31_5                                                                   (32'h1001abe4)
`define PV_REG_PCR_ENTRY_31_5                                                                       (32'hbe4)
`define CLP_PV_REG_PCR_ENTRY_31_6                                                                   (32'h1001abe8)
`define PV_REG_PCR_ENTRY_31_6                                                                       (32'hbe8)
`define CLP_PV_REG_PCR_ENTRY_31_7                                                                   (32'h1001abec)
`define PV_REG_PCR_ENTRY_31_7                                                                       (32'hbec)
`define CLP_PV_REG_PCR_ENTRY_31_8                                                                   (32'h1001abf0)
`define PV_REG_PCR_ENTRY_31_8                                                                       (32'hbf0)
`define CLP_PV_REG_PCR_ENTRY_31_9                                                                   (32'h1001abf4)
`define PV_REG_PCR_ENTRY_31_9                                                                       (32'hbf4)
`define CLP_PV_REG_PCR_ENTRY_31_10                                                                  (32'h1001abf8)
`define PV_REG_PCR_ENTRY_31_10                                                                      (32'hbf8)
`define CLP_PV_REG_PCR_ENTRY_31_11                                                                  (32'h1001abfc)
`define PV_REG_PCR_ENTRY_31_11                                                                      (32'hbfc)
`define CLP_DV_REG_BASE_ADDR                                                                        (32'h1001c000)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_0                                                            (32'h1001c000)
`define DV_REG_STICKYDATAVAULTCTRL_0                                                                (32'h0)
`define DV_REG_STICKYDATAVAULTCTRL_0_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_0_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_1                                                            (32'h1001c004)
`define DV_REG_STICKYDATAVAULTCTRL_1                                                                (32'h4)
`define DV_REG_STICKYDATAVAULTCTRL_1_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_1_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_2                                                            (32'h1001c008)
`define DV_REG_STICKYDATAVAULTCTRL_2                                                                (32'h8)
`define DV_REG_STICKYDATAVAULTCTRL_2_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_2_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_3                                                            (32'h1001c00c)
`define DV_REG_STICKYDATAVAULTCTRL_3                                                                (32'hc)
`define DV_REG_STICKYDATAVAULTCTRL_3_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_3_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_4                                                            (32'h1001c010)
`define DV_REG_STICKYDATAVAULTCTRL_4                                                                (32'h10)
`define DV_REG_STICKYDATAVAULTCTRL_4_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_4_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_5                                                            (32'h1001c014)
`define DV_REG_STICKYDATAVAULTCTRL_5                                                                (32'h14)
`define DV_REG_STICKYDATAVAULTCTRL_5_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_5_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_6                                                            (32'h1001c018)
`define DV_REG_STICKYDATAVAULTCTRL_6                                                                (32'h18)
`define DV_REG_STICKYDATAVAULTCTRL_6_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_6_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_7                                                            (32'h1001c01c)
`define DV_REG_STICKYDATAVAULTCTRL_7                                                                (32'h1c)
`define DV_REG_STICKYDATAVAULTCTRL_7_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_7_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_8                                                            (32'h1001c020)
`define DV_REG_STICKYDATAVAULTCTRL_8                                                                (32'h20)
`define DV_REG_STICKYDATAVAULTCTRL_8_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_8_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_9                                                            (32'h1001c024)
`define DV_REG_STICKYDATAVAULTCTRL_9                                                                (32'h24)
`define DV_REG_STICKYDATAVAULTCTRL_9_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_9_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_0                                                      (32'h1001c028)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_0                                                          (32'h28)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_1                                                      (32'h1001c02c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_1                                                          (32'h2c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_2                                                      (32'h1001c030)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_2                                                          (32'h30)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_3                                                      (32'h1001c034)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_3                                                          (32'h34)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_4                                                      (32'h1001c038)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_4                                                          (32'h38)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_5                                                      (32'h1001c03c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_5                                                          (32'h3c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_6                                                      (32'h1001c040)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_6                                                          (32'h40)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_7                                                      (32'h1001c044)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_7                                                          (32'h44)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_8                                                      (32'h1001c048)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_8                                                          (32'h48)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_9                                                      (32'h1001c04c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_9                                                          (32'h4c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_10                                                     (32'h1001c050)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_10                                                         (32'h50)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_11                                                     (32'h1001c054)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_11                                                         (32'h54)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_0                                                      (32'h1001c058)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_0                                                          (32'h58)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_1                                                      (32'h1001c05c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_1                                                          (32'h5c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_2                                                      (32'h1001c060)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_2                                                          (32'h60)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_3                                                      (32'h1001c064)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_3                                                          (32'h64)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_4                                                      (32'h1001c068)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_4                                                          (32'h68)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_5                                                      (32'h1001c06c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_5                                                          (32'h6c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_6                                                      (32'h1001c070)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_6                                                          (32'h70)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_7                                                      (32'h1001c074)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_7                                                          (32'h74)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_8                                                      (32'h1001c078)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_8                                                          (32'h78)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_9                                                      (32'h1001c07c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_9                                                          (32'h7c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_10                                                     (32'h1001c080)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_10                                                         (32'h80)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_11                                                     (32'h1001c084)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_11                                                         (32'h84)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_0                                                      (32'h1001c088)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_0                                                          (32'h88)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_1                                                      (32'h1001c08c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_1                                                          (32'h8c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_2                                                      (32'h1001c090)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_2                                                          (32'h90)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_3                                                      (32'h1001c094)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_3                                                          (32'h94)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_4                                                      (32'h1001c098)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_4                                                          (32'h98)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_5                                                      (32'h1001c09c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_5                                                          (32'h9c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_6                                                      (32'h1001c0a0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_6                                                          (32'ha0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_7                                                      (32'h1001c0a4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_7                                                          (32'ha4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_8                                                      (32'h1001c0a8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_8                                                          (32'ha8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_9                                                      (32'h1001c0ac)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_9                                                          (32'hac)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_10                                                     (32'h1001c0b0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_10                                                         (32'hb0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_11                                                     (32'h1001c0b4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_11                                                         (32'hb4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_0                                                      (32'h1001c0b8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_0                                                          (32'hb8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_1                                                      (32'h1001c0bc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_1                                                          (32'hbc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_2                                                      (32'h1001c0c0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_2                                                          (32'hc0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_3                                                      (32'h1001c0c4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_3                                                          (32'hc4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_4                                                      (32'h1001c0c8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_4                                                          (32'hc8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_5                                                      (32'h1001c0cc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_5                                                          (32'hcc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_6                                                      (32'h1001c0d0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_6                                                          (32'hd0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_7                                                      (32'h1001c0d4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_7                                                          (32'hd4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_8                                                      (32'h1001c0d8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_8                                                          (32'hd8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_9                                                      (32'h1001c0dc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_9                                                          (32'hdc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_10                                                     (32'h1001c0e0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_10                                                         (32'he0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_11                                                     (32'h1001c0e4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_11                                                         (32'he4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_0                                                      (32'h1001c0e8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_0                                                          (32'he8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_1                                                      (32'h1001c0ec)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_1                                                          (32'hec)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_2                                                      (32'h1001c0f0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_2                                                          (32'hf0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_3                                                      (32'h1001c0f4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_3                                                          (32'hf4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_4                                                      (32'h1001c0f8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_4                                                          (32'hf8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_5                                                      (32'h1001c0fc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_5                                                          (32'hfc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_6                                                      (32'h1001c100)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_6                                                          (32'h100)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_7                                                      (32'h1001c104)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_7                                                          (32'h104)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_8                                                      (32'h1001c108)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_8                                                          (32'h108)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_9                                                      (32'h1001c10c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_9                                                          (32'h10c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_10                                                     (32'h1001c110)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_10                                                         (32'h110)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_11                                                     (32'h1001c114)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_11                                                         (32'h114)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_0                                                      (32'h1001c118)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_0                                                          (32'h118)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_1                                                      (32'h1001c11c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_1                                                          (32'h11c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_2                                                      (32'h1001c120)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_2                                                          (32'h120)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_3                                                      (32'h1001c124)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_3                                                          (32'h124)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_4                                                      (32'h1001c128)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_4                                                          (32'h128)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_5                                                      (32'h1001c12c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_5                                                          (32'h12c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_6                                                      (32'h1001c130)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_6                                                          (32'h130)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_7                                                      (32'h1001c134)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_7                                                          (32'h134)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_8                                                      (32'h1001c138)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_8                                                          (32'h138)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_9                                                      (32'h1001c13c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_9                                                          (32'h13c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_10                                                     (32'h1001c140)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_10                                                         (32'h140)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_11                                                     (32'h1001c144)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_11                                                         (32'h144)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_0                                                      (32'h1001c148)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_0                                                          (32'h148)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_1                                                      (32'h1001c14c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_1                                                          (32'h14c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_2                                                      (32'h1001c150)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_2                                                          (32'h150)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_3                                                      (32'h1001c154)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_3                                                          (32'h154)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_4                                                      (32'h1001c158)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_4                                                          (32'h158)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_5                                                      (32'h1001c15c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_5                                                          (32'h15c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_6                                                      (32'h1001c160)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_6                                                          (32'h160)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_7                                                      (32'h1001c164)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_7                                                          (32'h164)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_8                                                      (32'h1001c168)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_8                                                          (32'h168)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_9                                                      (32'h1001c16c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_9                                                          (32'h16c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_10                                                     (32'h1001c170)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_10                                                         (32'h170)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_11                                                     (32'h1001c174)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_11                                                         (32'h174)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_0                                                      (32'h1001c178)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_0                                                          (32'h178)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_1                                                      (32'h1001c17c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_1                                                          (32'h17c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_2                                                      (32'h1001c180)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_2                                                          (32'h180)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_3                                                      (32'h1001c184)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_3                                                          (32'h184)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_4                                                      (32'h1001c188)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_4                                                          (32'h188)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_5                                                      (32'h1001c18c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_5                                                          (32'h18c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_6                                                      (32'h1001c190)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_6                                                          (32'h190)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_7                                                      (32'h1001c194)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_7                                                          (32'h194)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_8                                                      (32'h1001c198)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_8                                                          (32'h198)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_9                                                      (32'h1001c19c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_9                                                          (32'h19c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_10                                                     (32'h1001c1a0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_10                                                         (32'h1a0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_11                                                     (32'h1001c1a4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_11                                                         (32'h1a4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_0                                                      (32'h1001c1a8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_0                                                          (32'h1a8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_1                                                      (32'h1001c1ac)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_1                                                          (32'h1ac)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_2                                                      (32'h1001c1b0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_2                                                          (32'h1b0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_3                                                      (32'h1001c1b4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_3                                                          (32'h1b4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_4                                                      (32'h1001c1b8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_4                                                          (32'h1b8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_5                                                      (32'h1001c1bc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_5                                                          (32'h1bc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_6                                                      (32'h1001c1c0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_6                                                          (32'h1c0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_7                                                      (32'h1001c1c4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_7                                                          (32'h1c4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_8                                                      (32'h1001c1c8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_8                                                          (32'h1c8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_9                                                      (32'h1001c1cc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_9                                                          (32'h1cc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_10                                                     (32'h1001c1d0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_10                                                         (32'h1d0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_11                                                     (32'h1001c1d4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_11                                                         (32'h1d4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_0                                                      (32'h1001c1d8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_0                                                          (32'h1d8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_1                                                      (32'h1001c1dc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_1                                                          (32'h1dc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_2                                                      (32'h1001c1e0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_2                                                          (32'h1e0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_3                                                      (32'h1001c1e4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_3                                                          (32'h1e4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_4                                                      (32'h1001c1e8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_4                                                          (32'h1e8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_5                                                      (32'h1001c1ec)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_5                                                          (32'h1ec)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_6                                                      (32'h1001c1f0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_6                                                          (32'h1f0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_7                                                      (32'h1001c1f4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_7                                                          (32'h1f4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_8                                                      (32'h1001c1f8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_8                                                          (32'h1f8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_9                                                      (32'h1001c1fc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_9                                                          (32'h1fc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_10                                                     (32'h1001c200)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_10                                                         (32'h200)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_11                                                     (32'h1001c204)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_11                                                         (32'h204)
`define CLP_DV_REG_DATAVAULTCTRL_0                                                                  (32'h1001c208)
`define DV_REG_DATAVAULTCTRL_0                                                                      (32'h208)
`define DV_REG_DATAVAULTCTRL_0_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_0_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_1                                                                  (32'h1001c20c)
`define DV_REG_DATAVAULTCTRL_1                                                                      (32'h20c)
`define DV_REG_DATAVAULTCTRL_1_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_1_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_2                                                                  (32'h1001c210)
`define DV_REG_DATAVAULTCTRL_2                                                                      (32'h210)
`define DV_REG_DATAVAULTCTRL_2_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_2_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_3                                                                  (32'h1001c214)
`define DV_REG_DATAVAULTCTRL_3                                                                      (32'h214)
`define DV_REG_DATAVAULTCTRL_3_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_3_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_4                                                                  (32'h1001c218)
`define DV_REG_DATAVAULTCTRL_4                                                                      (32'h218)
`define DV_REG_DATAVAULTCTRL_4_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_4_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_5                                                                  (32'h1001c21c)
`define DV_REG_DATAVAULTCTRL_5                                                                      (32'h21c)
`define DV_REG_DATAVAULTCTRL_5_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_5_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_6                                                                  (32'h1001c220)
`define DV_REG_DATAVAULTCTRL_6                                                                      (32'h220)
`define DV_REG_DATAVAULTCTRL_6_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_6_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_7                                                                  (32'h1001c224)
`define DV_REG_DATAVAULTCTRL_7                                                                      (32'h224)
`define DV_REG_DATAVAULTCTRL_7_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_7_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_8                                                                  (32'h1001c228)
`define DV_REG_DATAVAULTCTRL_8                                                                      (32'h228)
`define DV_REG_DATAVAULTCTRL_8_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_8_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATAVAULTCTRL_9                                                                  (32'h1001c22c)
`define DV_REG_DATAVAULTCTRL_9                                                                      (32'h22c)
`define DV_REG_DATAVAULTCTRL_9_LOCK_ENTRY_LOW                                                       (0)
`define DV_REG_DATAVAULTCTRL_9_LOCK_ENTRY_MASK                                                      (32'h1)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_0                                                             (32'h1001c230)
`define DV_REG_DATA_VAULT_ENTRY_0_0                                                                 (32'h230)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_1                                                             (32'h1001c234)
`define DV_REG_DATA_VAULT_ENTRY_0_1                                                                 (32'h234)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_2                                                             (32'h1001c238)
`define DV_REG_DATA_VAULT_ENTRY_0_2                                                                 (32'h238)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_3                                                             (32'h1001c23c)
`define DV_REG_DATA_VAULT_ENTRY_0_3                                                                 (32'h23c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_4                                                             (32'h1001c240)
`define DV_REG_DATA_VAULT_ENTRY_0_4                                                                 (32'h240)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_5                                                             (32'h1001c244)
`define DV_REG_DATA_VAULT_ENTRY_0_5                                                                 (32'h244)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_6                                                             (32'h1001c248)
`define DV_REG_DATA_VAULT_ENTRY_0_6                                                                 (32'h248)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_7                                                             (32'h1001c24c)
`define DV_REG_DATA_VAULT_ENTRY_0_7                                                                 (32'h24c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_8                                                             (32'h1001c250)
`define DV_REG_DATA_VAULT_ENTRY_0_8                                                                 (32'h250)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_9                                                             (32'h1001c254)
`define DV_REG_DATA_VAULT_ENTRY_0_9                                                                 (32'h254)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_10                                                            (32'h1001c258)
`define DV_REG_DATA_VAULT_ENTRY_0_10                                                                (32'h258)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_11                                                            (32'h1001c25c)
`define DV_REG_DATA_VAULT_ENTRY_0_11                                                                (32'h25c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_0                                                             (32'h1001c260)
`define DV_REG_DATA_VAULT_ENTRY_1_0                                                                 (32'h260)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_1                                                             (32'h1001c264)
`define DV_REG_DATA_VAULT_ENTRY_1_1                                                                 (32'h264)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_2                                                             (32'h1001c268)
`define DV_REG_DATA_VAULT_ENTRY_1_2                                                                 (32'h268)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_3                                                             (32'h1001c26c)
`define DV_REG_DATA_VAULT_ENTRY_1_3                                                                 (32'h26c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_4                                                             (32'h1001c270)
`define DV_REG_DATA_VAULT_ENTRY_1_4                                                                 (32'h270)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_5                                                             (32'h1001c274)
`define DV_REG_DATA_VAULT_ENTRY_1_5                                                                 (32'h274)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_6                                                             (32'h1001c278)
`define DV_REG_DATA_VAULT_ENTRY_1_6                                                                 (32'h278)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_7                                                             (32'h1001c27c)
`define DV_REG_DATA_VAULT_ENTRY_1_7                                                                 (32'h27c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_8                                                             (32'h1001c280)
`define DV_REG_DATA_VAULT_ENTRY_1_8                                                                 (32'h280)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_9                                                             (32'h1001c284)
`define DV_REG_DATA_VAULT_ENTRY_1_9                                                                 (32'h284)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_10                                                            (32'h1001c288)
`define DV_REG_DATA_VAULT_ENTRY_1_10                                                                (32'h288)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_11                                                            (32'h1001c28c)
`define DV_REG_DATA_VAULT_ENTRY_1_11                                                                (32'h28c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_0                                                             (32'h1001c290)
`define DV_REG_DATA_VAULT_ENTRY_2_0                                                                 (32'h290)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_1                                                             (32'h1001c294)
`define DV_REG_DATA_VAULT_ENTRY_2_1                                                                 (32'h294)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_2                                                             (32'h1001c298)
`define DV_REG_DATA_VAULT_ENTRY_2_2                                                                 (32'h298)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_3                                                             (32'h1001c29c)
`define DV_REG_DATA_VAULT_ENTRY_2_3                                                                 (32'h29c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_4                                                             (32'h1001c2a0)
`define DV_REG_DATA_VAULT_ENTRY_2_4                                                                 (32'h2a0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_5                                                             (32'h1001c2a4)
`define DV_REG_DATA_VAULT_ENTRY_2_5                                                                 (32'h2a4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_6                                                             (32'h1001c2a8)
`define DV_REG_DATA_VAULT_ENTRY_2_6                                                                 (32'h2a8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_7                                                             (32'h1001c2ac)
`define DV_REG_DATA_VAULT_ENTRY_2_7                                                                 (32'h2ac)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_8                                                             (32'h1001c2b0)
`define DV_REG_DATA_VAULT_ENTRY_2_8                                                                 (32'h2b0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_9                                                             (32'h1001c2b4)
`define DV_REG_DATA_VAULT_ENTRY_2_9                                                                 (32'h2b4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_10                                                            (32'h1001c2b8)
`define DV_REG_DATA_VAULT_ENTRY_2_10                                                                (32'h2b8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_11                                                            (32'h1001c2bc)
`define DV_REG_DATA_VAULT_ENTRY_2_11                                                                (32'h2bc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_0                                                             (32'h1001c2c0)
`define DV_REG_DATA_VAULT_ENTRY_3_0                                                                 (32'h2c0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_1                                                             (32'h1001c2c4)
`define DV_REG_DATA_VAULT_ENTRY_3_1                                                                 (32'h2c4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_2                                                             (32'h1001c2c8)
`define DV_REG_DATA_VAULT_ENTRY_3_2                                                                 (32'h2c8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_3                                                             (32'h1001c2cc)
`define DV_REG_DATA_VAULT_ENTRY_3_3                                                                 (32'h2cc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_4                                                             (32'h1001c2d0)
`define DV_REG_DATA_VAULT_ENTRY_3_4                                                                 (32'h2d0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_5                                                             (32'h1001c2d4)
`define DV_REG_DATA_VAULT_ENTRY_3_5                                                                 (32'h2d4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_6                                                             (32'h1001c2d8)
`define DV_REG_DATA_VAULT_ENTRY_3_6                                                                 (32'h2d8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_7                                                             (32'h1001c2dc)
`define DV_REG_DATA_VAULT_ENTRY_3_7                                                                 (32'h2dc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_8                                                             (32'h1001c2e0)
`define DV_REG_DATA_VAULT_ENTRY_3_8                                                                 (32'h2e0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_9                                                             (32'h1001c2e4)
`define DV_REG_DATA_VAULT_ENTRY_3_9                                                                 (32'h2e4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_10                                                            (32'h1001c2e8)
`define DV_REG_DATA_VAULT_ENTRY_3_10                                                                (32'h2e8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_11                                                            (32'h1001c2ec)
`define DV_REG_DATA_VAULT_ENTRY_3_11                                                                (32'h2ec)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_0                                                             (32'h1001c2f0)
`define DV_REG_DATA_VAULT_ENTRY_4_0                                                                 (32'h2f0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_1                                                             (32'h1001c2f4)
`define DV_REG_DATA_VAULT_ENTRY_4_1                                                                 (32'h2f4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_2                                                             (32'h1001c2f8)
`define DV_REG_DATA_VAULT_ENTRY_4_2                                                                 (32'h2f8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_3                                                             (32'h1001c2fc)
`define DV_REG_DATA_VAULT_ENTRY_4_3                                                                 (32'h2fc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_4                                                             (32'h1001c300)
`define DV_REG_DATA_VAULT_ENTRY_4_4                                                                 (32'h300)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_5                                                             (32'h1001c304)
`define DV_REG_DATA_VAULT_ENTRY_4_5                                                                 (32'h304)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_6                                                             (32'h1001c308)
`define DV_REG_DATA_VAULT_ENTRY_4_6                                                                 (32'h308)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_7                                                             (32'h1001c30c)
`define DV_REG_DATA_VAULT_ENTRY_4_7                                                                 (32'h30c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_8                                                             (32'h1001c310)
`define DV_REG_DATA_VAULT_ENTRY_4_8                                                                 (32'h310)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_9                                                             (32'h1001c314)
`define DV_REG_DATA_VAULT_ENTRY_4_9                                                                 (32'h314)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_10                                                            (32'h1001c318)
`define DV_REG_DATA_VAULT_ENTRY_4_10                                                                (32'h318)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_11                                                            (32'h1001c31c)
`define DV_REG_DATA_VAULT_ENTRY_4_11                                                                (32'h31c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_0                                                             (32'h1001c320)
`define DV_REG_DATA_VAULT_ENTRY_5_0                                                                 (32'h320)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_1                                                             (32'h1001c324)
`define DV_REG_DATA_VAULT_ENTRY_5_1                                                                 (32'h324)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_2                                                             (32'h1001c328)
`define DV_REG_DATA_VAULT_ENTRY_5_2                                                                 (32'h328)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_3                                                             (32'h1001c32c)
`define DV_REG_DATA_VAULT_ENTRY_5_3                                                                 (32'h32c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_4                                                             (32'h1001c330)
`define DV_REG_DATA_VAULT_ENTRY_5_4                                                                 (32'h330)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_5                                                             (32'h1001c334)
`define DV_REG_DATA_VAULT_ENTRY_5_5                                                                 (32'h334)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_6                                                             (32'h1001c338)
`define DV_REG_DATA_VAULT_ENTRY_5_6                                                                 (32'h338)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_7                                                             (32'h1001c33c)
`define DV_REG_DATA_VAULT_ENTRY_5_7                                                                 (32'h33c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_8                                                             (32'h1001c340)
`define DV_REG_DATA_VAULT_ENTRY_5_8                                                                 (32'h340)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_9                                                             (32'h1001c344)
`define DV_REG_DATA_VAULT_ENTRY_5_9                                                                 (32'h344)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_10                                                            (32'h1001c348)
`define DV_REG_DATA_VAULT_ENTRY_5_10                                                                (32'h348)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_11                                                            (32'h1001c34c)
`define DV_REG_DATA_VAULT_ENTRY_5_11                                                                (32'h34c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_0                                                             (32'h1001c350)
`define DV_REG_DATA_VAULT_ENTRY_6_0                                                                 (32'h350)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_1                                                             (32'h1001c354)
`define DV_REG_DATA_VAULT_ENTRY_6_1                                                                 (32'h354)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_2                                                             (32'h1001c358)
`define DV_REG_DATA_VAULT_ENTRY_6_2                                                                 (32'h358)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_3                                                             (32'h1001c35c)
`define DV_REG_DATA_VAULT_ENTRY_6_3                                                                 (32'h35c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_4                                                             (32'h1001c360)
`define DV_REG_DATA_VAULT_ENTRY_6_4                                                                 (32'h360)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_5                                                             (32'h1001c364)
`define DV_REG_DATA_VAULT_ENTRY_6_5                                                                 (32'h364)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_6                                                             (32'h1001c368)
`define DV_REG_DATA_VAULT_ENTRY_6_6                                                                 (32'h368)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_7                                                             (32'h1001c36c)
`define DV_REG_DATA_VAULT_ENTRY_6_7                                                                 (32'h36c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_8                                                             (32'h1001c370)
`define DV_REG_DATA_VAULT_ENTRY_6_8                                                                 (32'h370)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_9                                                             (32'h1001c374)
`define DV_REG_DATA_VAULT_ENTRY_6_9                                                                 (32'h374)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_10                                                            (32'h1001c378)
`define DV_REG_DATA_VAULT_ENTRY_6_10                                                                (32'h378)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_11                                                            (32'h1001c37c)
`define DV_REG_DATA_VAULT_ENTRY_6_11                                                                (32'h37c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_0                                                             (32'h1001c380)
`define DV_REG_DATA_VAULT_ENTRY_7_0                                                                 (32'h380)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_1                                                             (32'h1001c384)
`define DV_REG_DATA_VAULT_ENTRY_7_1                                                                 (32'h384)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_2                                                             (32'h1001c388)
`define DV_REG_DATA_VAULT_ENTRY_7_2                                                                 (32'h388)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_3                                                             (32'h1001c38c)
`define DV_REG_DATA_VAULT_ENTRY_7_3                                                                 (32'h38c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_4                                                             (32'h1001c390)
`define DV_REG_DATA_VAULT_ENTRY_7_4                                                                 (32'h390)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_5                                                             (32'h1001c394)
`define DV_REG_DATA_VAULT_ENTRY_7_5                                                                 (32'h394)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_6                                                             (32'h1001c398)
`define DV_REG_DATA_VAULT_ENTRY_7_6                                                                 (32'h398)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_7                                                             (32'h1001c39c)
`define DV_REG_DATA_VAULT_ENTRY_7_7                                                                 (32'h39c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_8                                                             (32'h1001c3a0)
`define DV_REG_DATA_VAULT_ENTRY_7_8                                                                 (32'h3a0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_9                                                             (32'h1001c3a4)
`define DV_REG_DATA_VAULT_ENTRY_7_9                                                                 (32'h3a4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_10                                                            (32'h1001c3a8)
`define DV_REG_DATA_VAULT_ENTRY_7_10                                                                (32'h3a8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_11                                                            (32'h1001c3ac)
`define DV_REG_DATA_VAULT_ENTRY_7_11                                                                (32'h3ac)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_0                                                             (32'h1001c3b0)
`define DV_REG_DATA_VAULT_ENTRY_8_0                                                                 (32'h3b0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_1                                                             (32'h1001c3b4)
`define DV_REG_DATA_VAULT_ENTRY_8_1                                                                 (32'h3b4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_2                                                             (32'h1001c3b8)
`define DV_REG_DATA_VAULT_ENTRY_8_2                                                                 (32'h3b8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_3                                                             (32'h1001c3bc)
`define DV_REG_DATA_VAULT_ENTRY_8_3                                                                 (32'h3bc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_4                                                             (32'h1001c3c0)
`define DV_REG_DATA_VAULT_ENTRY_8_4                                                                 (32'h3c0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_5                                                             (32'h1001c3c4)
`define DV_REG_DATA_VAULT_ENTRY_8_5                                                                 (32'h3c4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_6                                                             (32'h1001c3c8)
`define DV_REG_DATA_VAULT_ENTRY_8_6                                                                 (32'h3c8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_7                                                             (32'h1001c3cc)
`define DV_REG_DATA_VAULT_ENTRY_8_7                                                                 (32'h3cc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_8                                                             (32'h1001c3d0)
`define DV_REG_DATA_VAULT_ENTRY_8_8                                                                 (32'h3d0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_9                                                             (32'h1001c3d4)
`define DV_REG_DATA_VAULT_ENTRY_8_9                                                                 (32'h3d4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_10                                                            (32'h1001c3d8)
`define DV_REG_DATA_VAULT_ENTRY_8_10                                                                (32'h3d8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_11                                                            (32'h1001c3dc)
`define DV_REG_DATA_VAULT_ENTRY_8_11                                                                (32'h3dc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_0                                                             (32'h1001c3e0)
`define DV_REG_DATA_VAULT_ENTRY_9_0                                                                 (32'h3e0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_1                                                             (32'h1001c3e4)
`define DV_REG_DATA_VAULT_ENTRY_9_1                                                                 (32'h3e4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_2                                                             (32'h1001c3e8)
`define DV_REG_DATA_VAULT_ENTRY_9_2                                                                 (32'h3e8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_3                                                             (32'h1001c3ec)
`define DV_REG_DATA_VAULT_ENTRY_9_3                                                                 (32'h3ec)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_4                                                             (32'h1001c3f0)
`define DV_REG_DATA_VAULT_ENTRY_9_4                                                                 (32'h3f0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_5                                                             (32'h1001c3f4)
`define DV_REG_DATA_VAULT_ENTRY_9_5                                                                 (32'h3f4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_6                                                             (32'h1001c3f8)
`define DV_REG_DATA_VAULT_ENTRY_9_6                                                                 (32'h3f8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_7                                                             (32'h1001c3fc)
`define DV_REG_DATA_VAULT_ENTRY_9_7                                                                 (32'h3fc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_8                                                             (32'h1001c400)
`define DV_REG_DATA_VAULT_ENTRY_9_8                                                                 (32'h400)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_9                                                             (32'h1001c404)
`define DV_REG_DATA_VAULT_ENTRY_9_9                                                                 (32'h404)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_10                                                            (32'h1001c408)
`define DV_REG_DATA_VAULT_ENTRY_9_10                                                                (32'h408)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_11                                                            (32'h1001c40c)
`define DV_REG_DATA_VAULT_ENTRY_9_11                                                                (32'h40c)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_0                                                         (32'h1001c410)
`define DV_REG_LOCKABLESCRATCHREGCTRL_0                                                             (32'h410)
`define DV_REG_LOCKABLESCRATCHREGCTRL_0_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_0_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_1                                                         (32'h1001c414)
`define DV_REG_LOCKABLESCRATCHREGCTRL_1                                                             (32'h414)
`define DV_REG_LOCKABLESCRATCHREGCTRL_1_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_1_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_2                                                         (32'h1001c418)
`define DV_REG_LOCKABLESCRATCHREGCTRL_2                                                             (32'h418)
`define DV_REG_LOCKABLESCRATCHREGCTRL_2_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_2_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_3                                                         (32'h1001c41c)
`define DV_REG_LOCKABLESCRATCHREGCTRL_3                                                             (32'h41c)
`define DV_REG_LOCKABLESCRATCHREGCTRL_3_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_3_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_4                                                         (32'h1001c420)
`define DV_REG_LOCKABLESCRATCHREGCTRL_4                                                             (32'h420)
`define DV_REG_LOCKABLESCRATCHREGCTRL_4_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_4_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_5                                                         (32'h1001c424)
`define DV_REG_LOCKABLESCRATCHREGCTRL_5                                                             (32'h424)
`define DV_REG_LOCKABLESCRATCHREGCTRL_5_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_5_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_6                                                         (32'h1001c428)
`define DV_REG_LOCKABLESCRATCHREGCTRL_6                                                             (32'h428)
`define DV_REG_LOCKABLESCRATCHREGCTRL_6_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_6_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_7                                                         (32'h1001c42c)
`define DV_REG_LOCKABLESCRATCHREGCTRL_7                                                             (32'h42c)
`define DV_REG_LOCKABLESCRATCHREGCTRL_7_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_7_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_8                                                         (32'h1001c430)
`define DV_REG_LOCKABLESCRATCHREGCTRL_8                                                             (32'h430)
`define DV_REG_LOCKABLESCRATCHREGCTRL_8_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_8_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_9                                                         (32'h1001c434)
`define DV_REG_LOCKABLESCRATCHREGCTRL_9                                                             (32'h434)
`define DV_REG_LOCKABLESCRATCHREGCTRL_9_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_LOCKABLESCRATCHREGCTRL_9_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_LOCKABLESCRATCHREG_0                                                             (32'h1001c438)
`define DV_REG_LOCKABLESCRATCHREG_0                                                                 (32'h438)
`define CLP_DV_REG_LOCKABLESCRATCHREG_1                                                             (32'h1001c43c)
`define DV_REG_LOCKABLESCRATCHREG_1                                                                 (32'h43c)
`define CLP_DV_REG_LOCKABLESCRATCHREG_2                                                             (32'h1001c440)
`define DV_REG_LOCKABLESCRATCHREG_2                                                                 (32'h440)
`define CLP_DV_REG_LOCKABLESCRATCHREG_3                                                             (32'h1001c444)
`define DV_REG_LOCKABLESCRATCHREG_3                                                                 (32'h444)
`define CLP_DV_REG_LOCKABLESCRATCHREG_4                                                             (32'h1001c448)
`define DV_REG_LOCKABLESCRATCHREG_4                                                                 (32'h448)
`define CLP_DV_REG_LOCKABLESCRATCHREG_5                                                             (32'h1001c44c)
`define DV_REG_LOCKABLESCRATCHREG_5                                                                 (32'h44c)
`define CLP_DV_REG_LOCKABLESCRATCHREG_6                                                             (32'h1001c450)
`define DV_REG_LOCKABLESCRATCHREG_6                                                                 (32'h450)
`define CLP_DV_REG_LOCKABLESCRATCHREG_7                                                             (32'h1001c454)
`define DV_REG_LOCKABLESCRATCHREG_7                                                                 (32'h454)
`define CLP_DV_REG_LOCKABLESCRATCHREG_8                                                             (32'h1001c458)
`define DV_REG_LOCKABLESCRATCHREG_8                                                                 (32'h458)
`define CLP_DV_REG_LOCKABLESCRATCHREG_9                                                             (32'h1001c45c)
`define DV_REG_LOCKABLESCRATCHREG_9                                                                 (32'h45c)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_0                                                     (32'h1001c460)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_0                                                         (32'h460)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_1                                                     (32'h1001c464)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_1                                                         (32'h464)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_2                                                     (32'h1001c468)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_2                                                         (32'h468)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_3                                                     (32'h1001c46c)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_3                                                         (32'h46c)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_4                                                     (32'h1001c470)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_4                                                         (32'h470)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_5                                                     (32'h1001c474)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_5                                                         (32'h474)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_6                                                     (32'h1001c478)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_6                                                         (32'h478)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_7                                                     (32'h1001c47c)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_7                                                         (32'h47c)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0                                                   (32'h1001c480)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0                                                       (32'h480)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1                                                   (32'h1001c484)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1                                                       (32'h484)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2                                                   (32'h1001c488)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2                                                       (32'h488)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3                                                   (32'h1001c48c)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3                                                       (32'h48c)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4                                                   (32'h1001c490)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4                                                       (32'h490)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5                                                   (32'h1001c494)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5                                                       (32'h494)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6                                                   (32'h1001c498)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6                                                       (32'h498)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7                                                   (32'h1001c49c)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7                                                       (32'h49c)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_0                                                       (32'h1001c4a0)
`define DV_REG_STICKYLOCKABLESCRATCHREG_0                                                           (32'h4a0)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_1                                                       (32'h1001c4a4)
`define DV_REG_STICKYLOCKABLESCRATCHREG_1                                                           (32'h4a4)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_2                                                       (32'h1001c4a8)
`define DV_REG_STICKYLOCKABLESCRATCHREG_2                                                           (32'h4a8)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_3                                                       (32'h1001c4ac)
`define DV_REG_STICKYLOCKABLESCRATCHREG_3                                                           (32'h4ac)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_4                                                       (32'h1001c4b0)
`define DV_REG_STICKYLOCKABLESCRATCHREG_4                                                           (32'h4b0)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_5                                                       (32'h1001c4b4)
`define DV_REG_STICKYLOCKABLESCRATCHREG_5                                                           (32'h4b4)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_6                                                       (32'h1001c4b8)
`define DV_REG_STICKYLOCKABLESCRATCHREG_6                                                           (32'h4b8)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_7                                                       (32'h1001c4bc)
`define DV_REG_STICKYLOCKABLESCRATCHREG_7                                                           (32'h4bc)
`define CLP_SHA512_REG_BASE_ADDR                                                                    (32'h10020000)
`define CLP_SHA512_REG_SHA512_NAME_0                                                                (32'h10020000)
`define SHA512_REG_SHA512_NAME_0                                                                    (32'h0)
`define CLP_SHA512_REG_SHA512_NAME_1                                                                (32'h10020004)
`define SHA512_REG_SHA512_NAME_1                                                                    (32'h4)
`define CLP_SHA512_REG_SHA512_VERSION_0                                                             (32'h10020008)
`define SHA512_REG_SHA512_VERSION_0                                                                 (32'h8)
`define CLP_SHA512_REG_SHA512_VERSION_1                                                             (32'h1002000c)
`define SHA512_REG_SHA512_VERSION_1                                                                 (32'hc)
`define CLP_SHA512_REG_SHA512_CTRL                                                                  (32'h10020010)
`define SHA512_REG_SHA512_CTRL                                                                      (32'h10)
`define SHA512_REG_SHA512_CTRL_INIT_LOW                                                             (0)
`define SHA512_REG_SHA512_CTRL_INIT_MASK                                                            (32'h1)
`define SHA512_REG_SHA512_CTRL_NEXT_LOW                                                             (1)
`define SHA512_REG_SHA512_CTRL_NEXT_MASK                                                            (32'h2)
`define SHA512_REG_SHA512_CTRL_MODE_LOW                                                             (2)
`define SHA512_REG_SHA512_CTRL_MODE_MASK                                                            (32'hc)
`define SHA512_REG_SHA512_CTRL_ZEROIZE_LOW                                                          (4)
`define SHA512_REG_SHA512_CTRL_ZEROIZE_MASK                                                         (32'h10)
`define SHA512_REG_SHA512_CTRL_LAST_LOW                                                             (5)
`define SHA512_REG_SHA512_CTRL_LAST_MASK                                                            (32'h20)
`define CLP_SHA512_REG_SHA512_STATUS                                                                (32'h10020018)
`define SHA512_REG_SHA512_STATUS                                                                    (32'h18)
`define SHA512_REG_SHA512_STATUS_READY_LOW                                                          (0)
`define SHA512_REG_SHA512_STATUS_READY_MASK                                                         (32'h1)
`define SHA512_REG_SHA512_STATUS_VALID_LOW                                                          (1)
`define SHA512_REG_SHA512_STATUS_VALID_MASK                                                         (32'h2)
`define CLP_SHA512_REG_SHA512_BLOCK_0                                                               (32'h10020080)
`define SHA512_REG_SHA512_BLOCK_0                                                                   (32'h80)
`define CLP_SHA512_REG_SHA512_BLOCK_1                                                               (32'h10020084)
`define SHA512_REG_SHA512_BLOCK_1                                                                   (32'h84)
`define CLP_SHA512_REG_SHA512_BLOCK_2                                                               (32'h10020088)
`define SHA512_REG_SHA512_BLOCK_2                                                                   (32'h88)
`define CLP_SHA512_REG_SHA512_BLOCK_3                                                               (32'h1002008c)
`define SHA512_REG_SHA512_BLOCK_3                                                                   (32'h8c)
`define CLP_SHA512_REG_SHA512_BLOCK_4                                                               (32'h10020090)
`define SHA512_REG_SHA512_BLOCK_4                                                                   (32'h90)
`define CLP_SHA512_REG_SHA512_BLOCK_5                                                               (32'h10020094)
`define SHA512_REG_SHA512_BLOCK_5                                                                   (32'h94)
`define CLP_SHA512_REG_SHA512_BLOCK_6                                                               (32'h10020098)
`define SHA512_REG_SHA512_BLOCK_6                                                                   (32'h98)
`define CLP_SHA512_REG_SHA512_BLOCK_7                                                               (32'h1002009c)
`define SHA512_REG_SHA512_BLOCK_7                                                                   (32'h9c)
`define CLP_SHA512_REG_SHA512_BLOCK_8                                                               (32'h100200a0)
`define SHA512_REG_SHA512_BLOCK_8                                                                   (32'ha0)
`define CLP_SHA512_REG_SHA512_BLOCK_9                                                               (32'h100200a4)
`define SHA512_REG_SHA512_BLOCK_9                                                                   (32'ha4)
`define CLP_SHA512_REG_SHA512_BLOCK_10                                                              (32'h100200a8)
`define SHA512_REG_SHA512_BLOCK_10                                                                  (32'ha8)
`define CLP_SHA512_REG_SHA512_BLOCK_11                                                              (32'h100200ac)
`define SHA512_REG_SHA512_BLOCK_11                                                                  (32'hac)
`define CLP_SHA512_REG_SHA512_BLOCK_12                                                              (32'h100200b0)
`define SHA512_REG_SHA512_BLOCK_12                                                                  (32'hb0)
`define CLP_SHA512_REG_SHA512_BLOCK_13                                                              (32'h100200b4)
`define SHA512_REG_SHA512_BLOCK_13                                                                  (32'hb4)
`define CLP_SHA512_REG_SHA512_BLOCK_14                                                              (32'h100200b8)
`define SHA512_REG_SHA512_BLOCK_14                                                                  (32'hb8)
`define CLP_SHA512_REG_SHA512_BLOCK_15                                                              (32'h100200bc)
`define SHA512_REG_SHA512_BLOCK_15                                                                  (32'hbc)
`define CLP_SHA512_REG_SHA512_BLOCK_16                                                              (32'h100200c0)
`define SHA512_REG_SHA512_BLOCK_16                                                                  (32'hc0)
`define CLP_SHA512_REG_SHA512_BLOCK_17                                                              (32'h100200c4)
`define SHA512_REG_SHA512_BLOCK_17                                                                  (32'hc4)
`define CLP_SHA512_REG_SHA512_BLOCK_18                                                              (32'h100200c8)
`define SHA512_REG_SHA512_BLOCK_18                                                                  (32'hc8)
`define CLP_SHA512_REG_SHA512_BLOCK_19                                                              (32'h100200cc)
`define SHA512_REG_SHA512_BLOCK_19                                                                  (32'hcc)
`define CLP_SHA512_REG_SHA512_BLOCK_20                                                              (32'h100200d0)
`define SHA512_REG_SHA512_BLOCK_20                                                                  (32'hd0)
`define CLP_SHA512_REG_SHA512_BLOCK_21                                                              (32'h100200d4)
`define SHA512_REG_SHA512_BLOCK_21                                                                  (32'hd4)
`define CLP_SHA512_REG_SHA512_BLOCK_22                                                              (32'h100200d8)
`define SHA512_REG_SHA512_BLOCK_22                                                                  (32'hd8)
`define CLP_SHA512_REG_SHA512_BLOCK_23                                                              (32'h100200dc)
`define SHA512_REG_SHA512_BLOCK_23                                                                  (32'hdc)
`define CLP_SHA512_REG_SHA512_BLOCK_24                                                              (32'h100200e0)
`define SHA512_REG_SHA512_BLOCK_24                                                                  (32'he0)
`define CLP_SHA512_REG_SHA512_BLOCK_25                                                              (32'h100200e4)
`define SHA512_REG_SHA512_BLOCK_25                                                                  (32'he4)
`define CLP_SHA512_REG_SHA512_BLOCK_26                                                              (32'h100200e8)
`define SHA512_REG_SHA512_BLOCK_26                                                                  (32'he8)
`define CLP_SHA512_REG_SHA512_BLOCK_27                                                              (32'h100200ec)
`define SHA512_REG_SHA512_BLOCK_27                                                                  (32'hec)
`define CLP_SHA512_REG_SHA512_BLOCK_28                                                              (32'h100200f0)
`define SHA512_REG_SHA512_BLOCK_28                                                                  (32'hf0)
`define CLP_SHA512_REG_SHA512_BLOCK_29                                                              (32'h100200f4)
`define SHA512_REG_SHA512_BLOCK_29                                                                  (32'hf4)
`define CLP_SHA512_REG_SHA512_BLOCK_30                                                              (32'h100200f8)
`define SHA512_REG_SHA512_BLOCK_30                                                                  (32'hf8)
`define CLP_SHA512_REG_SHA512_BLOCK_31                                                              (32'h100200fc)
`define SHA512_REG_SHA512_BLOCK_31                                                                  (32'hfc)
`define CLP_SHA512_REG_SHA512_DIGEST_0                                                              (32'h10020100)
`define SHA512_REG_SHA512_DIGEST_0                                                                  (32'h100)
`define CLP_SHA512_REG_SHA512_DIGEST_1                                                              (32'h10020104)
`define SHA512_REG_SHA512_DIGEST_1                                                                  (32'h104)
`define CLP_SHA512_REG_SHA512_DIGEST_2                                                              (32'h10020108)
`define SHA512_REG_SHA512_DIGEST_2                                                                  (32'h108)
`define CLP_SHA512_REG_SHA512_DIGEST_3                                                              (32'h1002010c)
`define SHA512_REG_SHA512_DIGEST_3                                                                  (32'h10c)
`define CLP_SHA512_REG_SHA512_DIGEST_4                                                              (32'h10020110)
`define SHA512_REG_SHA512_DIGEST_4                                                                  (32'h110)
`define CLP_SHA512_REG_SHA512_DIGEST_5                                                              (32'h10020114)
`define SHA512_REG_SHA512_DIGEST_5                                                                  (32'h114)
`define CLP_SHA512_REG_SHA512_DIGEST_6                                                              (32'h10020118)
`define SHA512_REG_SHA512_DIGEST_6                                                                  (32'h118)
`define CLP_SHA512_REG_SHA512_DIGEST_7                                                              (32'h1002011c)
`define SHA512_REG_SHA512_DIGEST_7                                                                  (32'h11c)
`define CLP_SHA512_REG_SHA512_DIGEST_8                                                              (32'h10020120)
`define SHA512_REG_SHA512_DIGEST_8                                                                  (32'h120)
`define CLP_SHA512_REG_SHA512_DIGEST_9                                                              (32'h10020124)
`define SHA512_REG_SHA512_DIGEST_9                                                                  (32'h124)
`define CLP_SHA512_REG_SHA512_DIGEST_10                                                             (32'h10020128)
`define SHA512_REG_SHA512_DIGEST_10                                                                 (32'h128)
`define CLP_SHA512_REG_SHA512_DIGEST_11                                                             (32'h1002012c)
`define SHA512_REG_SHA512_DIGEST_11                                                                 (32'h12c)
`define CLP_SHA512_REG_SHA512_DIGEST_12                                                             (32'h10020130)
`define SHA512_REG_SHA512_DIGEST_12                                                                 (32'h130)
`define CLP_SHA512_REG_SHA512_DIGEST_13                                                             (32'h10020134)
`define SHA512_REG_SHA512_DIGEST_13                                                                 (32'h134)
`define CLP_SHA512_REG_SHA512_DIGEST_14                                                             (32'h10020138)
`define SHA512_REG_SHA512_DIGEST_14                                                                 (32'h138)
`define CLP_SHA512_REG_SHA512_DIGEST_15                                                             (32'h1002013c)
`define SHA512_REG_SHA512_DIGEST_15                                                                 (32'h13c)
`define CLP_SHA512_REG_SHA512_VAULT_RD_CTRL                                                         (32'h10020600)
`define SHA512_REG_SHA512_VAULT_RD_CTRL                                                             (32'h600)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_READ_EN_LOW                                                 (0)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_READ_EN_MASK                                                (32'h1)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_READ_ENTRY_LOW                                              (1)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_READ_ENTRY_MASK                                             (32'h3e)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_PCR_HASH_EXTEND_LOW                                         (6)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_PCR_HASH_EXTEND_MASK                                        (32'h40)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_RSVD_LOW                                                    (7)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_RSVD_MASK                                                   (32'hffffff80)
`define CLP_SHA512_REG_SHA512_VAULT_RD_STATUS                                                       (32'h10020604)
`define SHA512_REG_SHA512_VAULT_RD_STATUS                                                           (32'h604)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_READY_LOW                                                 (0)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_READY_MASK                                                (32'h1)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_VALID_LOW                                                 (1)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_VALID_MASK                                                (32'h2)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_ERROR_LOW                                                 (2)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_ERROR_MASK                                                (32'h3fc)
`define CLP_SHA512_REG_SHA512_KV_WR_CTRL                                                            (32'h10020608)
`define SHA512_REG_SHA512_KV_WR_CTRL                                                                (32'h608)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_EN_LOW                                                   (0)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_EN_MASK                                                  (32'h1)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_ENTRY_LOW                                                (1)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_ENTRY_MASK                                               (32'h3e)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_KEY_DEST_VALID_LOW                                        (6)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_KEY_DEST_VALID_MASK                                       (32'h40)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                      (7)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                     (32'h80)
`define SHA512_REG_SHA512_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_LOW                                       (8)
`define SHA512_REG_SHA512_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_MASK                                      (32'h100)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_PKEY_DEST_VALID_LOW                                        (9)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_PKEY_DEST_VALID_MASK                                       (32'h200)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_SEED_DEST_VALID_LOW                                        (10)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_SEED_DEST_VALID_MASK                                       (32'h400)
`define SHA512_REG_SHA512_KV_WR_CTRL_RSVD_LOW                                                       (11)
`define SHA512_REG_SHA512_KV_WR_CTRL_RSVD_MASK                                                      (32'hfffff800)
`define CLP_SHA512_REG_SHA512_KV_WR_STATUS                                                          (32'h1002060c)
`define SHA512_REG_SHA512_KV_WR_STATUS                                                              (32'h60c)
`define SHA512_REG_SHA512_KV_WR_STATUS_READY_LOW                                                    (0)
`define SHA512_REG_SHA512_KV_WR_STATUS_READY_MASK                                                   (32'h1)
`define SHA512_REG_SHA512_KV_WR_STATUS_VALID_LOW                                                    (1)
`define SHA512_REG_SHA512_KV_WR_STATUS_VALID_MASK                                                   (32'h2)
`define SHA512_REG_SHA512_KV_WR_STATUS_ERROR_LOW                                                    (2)
`define SHA512_REG_SHA512_KV_WR_STATUS_ERROR_MASK                                                   (32'h3fc)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_0                                                  (32'h10020610)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_0                                                      (32'h610)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_1                                                  (32'h10020614)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_1                                                      (32'h614)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_2                                                  (32'h10020618)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_2                                                      (32'h618)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_3                                                  (32'h1002061c)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_3                                                      (32'h61c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_4                                                  (32'h10020620)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_4                                                      (32'h620)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_5                                                  (32'h10020624)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_5                                                      (32'h624)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_6                                                  (32'h10020628)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_6                                                      (32'h628)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_7                                                  (32'h1002062c)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_7                                                      (32'h62c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_CTRL                                                     (32'h10020630)
`define SHA512_REG_SHA512_GEN_PCR_HASH_CTRL                                                         (32'h630)
`define SHA512_REG_SHA512_GEN_PCR_HASH_CTRL_START_LOW                                               (0)
`define SHA512_REG_SHA512_GEN_PCR_HASH_CTRL_START_MASK                                              (32'h1)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_STATUS                                                   (32'h10020634)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS                                                       (32'h634)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS_READY_LOW                                             (0)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS_READY_MASK                                            (32'h1)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS_VALID_LOW                                             (1)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS_VALID_MASK                                            (32'h2)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_0                                                 (32'h10020638)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_0                                                     (32'h638)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_1                                                 (32'h1002063c)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_1                                                     (32'h63c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_2                                                 (32'h10020640)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_2                                                     (32'h640)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_3                                                 (32'h10020644)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_3                                                     (32'h644)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_4                                                 (32'h10020648)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_4                                                     (32'h648)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_5                                                 (32'h1002064c)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_5                                                     (32'h64c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_6                                                 (32'h10020650)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_6                                                     (32'h650)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_7                                                 (32'h10020654)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_7                                                     (32'h654)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_8                                                 (32'h10020658)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_8                                                     (32'h658)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_9                                                 (32'h1002065c)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_9                                                     (32'h65c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_10                                                (32'h10020660)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_10                                                    (32'h660)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_11                                                (32'h10020664)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_11                                                    (32'h664)
`define CLP_SHA512_REG_INTR_BLOCK_RF_START                                                          (32'h10020800)
`define CLP_SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h10020800)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                   (32'h800)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                      (0)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                     (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                      (1)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                     (32'h2)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h10020804)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                    (32'h804)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                      (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                     (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                      (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                     (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                      (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                     (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                      (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                     (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h10020808)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                    (32'h808)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                              (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                             (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h1002080c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                (32'h80c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h10020810)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                (32'h810)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h10020814)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                              (32'h814)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                               (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                              (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                               (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                              (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                               (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                              (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                               (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                              (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h10020818)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                              (32'h818)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                       (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                      (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h1002081c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                  (32'h81c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                  (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                 (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                  (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                 (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                  (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                 (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                  (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                 (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h10020820)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                  (32'h820)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                          (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                         (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h10020900)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                (32'h900)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h10020904)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                (32'h904)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h10020908)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                (32'h908)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h1002090c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                (32'h90c)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h10020980)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                        (32'h980)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'h10020a00)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                           (32'ha00)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'h10020a04)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                           (32'ha04)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'h10020a08)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                           (32'ha08)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'h10020a0c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                           (32'ha0c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'h10020a10)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                   (32'ha10)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_SHA256_REG_BASE_ADDR                                                                    (32'h10028000)
`define CLP_SHA256_REG_SHA256_NAME_0                                                                (32'h10028000)
`define SHA256_REG_SHA256_NAME_0                                                                    (32'h0)
`define CLP_SHA256_REG_SHA256_NAME_1                                                                (32'h10028004)
`define SHA256_REG_SHA256_NAME_1                                                                    (32'h4)
`define CLP_SHA256_REG_SHA256_VERSION_0                                                             (32'h10028008)
`define SHA256_REG_SHA256_VERSION_0                                                                 (32'h8)
`define CLP_SHA256_REG_SHA256_VERSION_1                                                             (32'h1002800c)
`define SHA256_REG_SHA256_VERSION_1                                                                 (32'hc)
`define CLP_SHA256_REG_SHA256_CTRL                                                                  (32'h10028010)
`define SHA256_REG_SHA256_CTRL                                                                      (32'h10)
`define SHA256_REG_SHA256_CTRL_INIT_LOW                                                             (0)
`define SHA256_REG_SHA256_CTRL_INIT_MASK                                                            (32'h1)
`define SHA256_REG_SHA256_CTRL_NEXT_LOW                                                             (1)
`define SHA256_REG_SHA256_CTRL_NEXT_MASK                                                            (32'h2)
`define SHA256_REG_SHA256_CTRL_MODE_LOW                                                             (2)
`define SHA256_REG_SHA256_CTRL_MODE_MASK                                                            (32'h4)
`define SHA256_REG_SHA256_CTRL_ZEROIZE_LOW                                                          (3)
`define SHA256_REG_SHA256_CTRL_ZEROIZE_MASK                                                         (32'h8)
`define SHA256_REG_SHA256_CTRL_WNTZ_MODE_LOW                                                        (4)
`define SHA256_REG_SHA256_CTRL_WNTZ_MODE_MASK                                                       (32'h10)
`define SHA256_REG_SHA256_CTRL_WNTZ_W_LOW                                                           (5)
`define SHA256_REG_SHA256_CTRL_WNTZ_W_MASK                                                          (32'h1e0)
`define SHA256_REG_SHA256_CTRL_WNTZ_N_MODE_LOW                                                      (9)
`define SHA256_REG_SHA256_CTRL_WNTZ_N_MODE_MASK                                                     (32'h200)
`define CLP_SHA256_REG_SHA256_STATUS                                                                (32'h10028018)
`define SHA256_REG_SHA256_STATUS                                                                    (32'h18)
`define SHA256_REG_SHA256_STATUS_READY_LOW                                                          (0)
`define SHA256_REG_SHA256_STATUS_READY_MASK                                                         (32'h1)
`define SHA256_REG_SHA256_STATUS_VALID_LOW                                                          (1)
`define SHA256_REG_SHA256_STATUS_VALID_MASK                                                         (32'h2)
`define SHA256_REG_SHA256_STATUS_WNTZ_BUSY_LOW                                                      (2)
`define SHA256_REG_SHA256_STATUS_WNTZ_BUSY_MASK                                                     (32'h4)
`define CLP_SHA256_REG_SHA256_BLOCK_0                                                               (32'h10028080)
`define SHA256_REG_SHA256_BLOCK_0                                                                   (32'h80)
`define CLP_SHA256_REG_SHA256_BLOCK_1                                                               (32'h10028084)
`define SHA256_REG_SHA256_BLOCK_1                                                                   (32'h84)
`define CLP_SHA256_REG_SHA256_BLOCK_2                                                               (32'h10028088)
`define SHA256_REG_SHA256_BLOCK_2                                                                   (32'h88)
`define CLP_SHA256_REG_SHA256_BLOCK_3                                                               (32'h1002808c)
`define SHA256_REG_SHA256_BLOCK_3                                                                   (32'h8c)
`define CLP_SHA256_REG_SHA256_BLOCK_4                                                               (32'h10028090)
`define SHA256_REG_SHA256_BLOCK_4                                                                   (32'h90)
`define CLP_SHA256_REG_SHA256_BLOCK_5                                                               (32'h10028094)
`define SHA256_REG_SHA256_BLOCK_5                                                                   (32'h94)
`define CLP_SHA256_REG_SHA256_BLOCK_6                                                               (32'h10028098)
`define SHA256_REG_SHA256_BLOCK_6                                                                   (32'h98)
`define CLP_SHA256_REG_SHA256_BLOCK_7                                                               (32'h1002809c)
`define SHA256_REG_SHA256_BLOCK_7                                                                   (32'h9c)
`define CLP_SHA256_REG_SHA256_BLOCK_8                                                               (32'h100280a0)
`define SHA256_REG_SHA256_BLOCK_8                                                                   (32'ha0)
`define CLP_SHA256_REG_SHA256_BLOCK_9                                                               (32'h100280a4)
`define SHA256_REG_SHA256_BLOCK_9                                                                   (32'ha4)
`define CLP_SHA256_REG_SHA256_BLOCK_10                                                              (32'h100280a8)
`define SHA256_REG_SHA256_BLOCK_10                                                                  (32'ha8)
`define CLP_SHA256_REG_SHA256_BLOCK_11                                                              (32'h100280ac)
`define SHA256_REG_SHA256_BLOCK_11                                                                  (32'hac)
`define CLP_SHA256_REG_SHA256_BLOCK_12                                                              (32'h100280b0)
`define SHA256_REG_SHA256_BLOCK_12                                                                  (32'hb0)
`define CLP_SHA256_REG_SHA256_BLOCK_13                                                              (32'h100280b4)
`define SHA256_REG_SHA256_BLOCK_13                                                                  (32'hb4)
`define CLP_SHA256_REG_SHA256_BLOCK_14                                                              (32'h100280b8)
`define SHA256_REG_SHA256_BLOCK_14                                                                  (32'hb8)
`define CLP_SHA256_REG_SHA256_BLOCK_15                                                              (32'h100280bc)
`define SHA256_REG_SHA256_BLOCK_15                                                                  (32'hbc)
`define CLP_SHA256_REG_SHA256_DIGEST_0                                                              (32'h10028100)
`define SHA256_REG_SHA256_DIGEST_0                                                                  (32'h100)
`define CLP_SHA256_REG_SHA256_DIGEST_1                                                              (32'h10028104)
`define SHA256_REG_SHA256_DIGEST_1                                                                  (32'h104)
`define CLP_SHA256_REG_SHA256_DIGEST_2                                                              (32'h10028108)
`define SHA256_REG_SHA256_DIGEST_2                                                                  (32'h108)
`define CLP_SHA256_REG_SHA256_DIGEST_3                                                              (32'h1002810c)
`define SHA256_REG_SHA256_DIGEST_3                                                                  (32'h10c)
`define CLP_SHA256_REG_SHA256_DIGEST_4                                                              (32'h10028110)
`define SHA256_REG_SHA256_DIGEST_4                                                                  (32'h110)
`define CLP_SHA256_REG_SHA256_DIGEST_5                                                              (32'h10028114)
`define SHA256_REG_SHA256_DIGEST_5                                                                  (32'h114)
`define CLP_SHA256_REG_SHA256_DIGEST_6                                                              (32'h10028118)
`define SHA256_REG_SHA256_DIGEST_6                                                                  (32'h118)
`define CLP_SHA256_REG_SHA256_DIGEST_7                                                              (32'h1002811c)
`define SHA256_REG_SHA256_DIGEST_7                                                                  (32'h11c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_START                                                          (32'h10028800)
`define CLP_SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h10028800)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                   (32'h800)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                      (0)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                     (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                      (1)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                     (32'h2)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h10028804)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                    (32'h804)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                      (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                     (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                      (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                     (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                      (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                     (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                      (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                     (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h10028808)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                    (32'h808)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                              (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                             (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h1002880c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                (32'h80c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h10028810)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                (32'h810)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h10028814)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                              (32'h814)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                               (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                              (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                               (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                              (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                               (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                              (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                               (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                              (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h10028818)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                              (32'h818)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                       (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                      (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h1002881c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                  (32'h81c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                  (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                 (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                  (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                 (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                  (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                 (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                  (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                 (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h10028820)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                  (32'h820)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                          (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                         (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h10028900)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                (32'h900)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h10028904)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                (32'h904)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h10028908)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                (32'h908)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h1002890c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                (32'h90c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h10028980)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                        (32'h980)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'h10028a00)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                           (32'ha00)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'h10028a04)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                           (32'ha04)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'h10028a08)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                           (32'ha08)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'h10028a0c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                           (32'ha0c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'h10028a10)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                   (32'ha10)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_MLDSA_REG_BASE_ADDR                                                                     (32'h10030000)
`define CLP_MLDSA_REG_MLDSA_NAME_0                                                                  (32'h10030000)
`define MLDSA_REG_MLDSA_NAME_0                                                                      (32'h0)
`define CLP_MLDSA_REG_MLDSA_NAME_1                                                                  (32'h10030004)
`define MLDSA_REG_MLDSA_NAME_1                                                                      (32'h4)
`define CLP_MLDSA_REG_MLDSA_VERSION_0                                                               (32'h10030008)
`define MLDSA_REG_MLDSA_VERSION_0                                                                   (32'h8)
`define CLP_MLDSA_REG_MLDSA_VERSION_1                                                               (32'h1003000c)
`define MLDSA_REG_MLDSA_VERSION_1                                                                   (32'hc)
`define CLP_MLDSA_REG_MLDSA_CTRL                                                                    (32'h10030010)
`define MLDSA_REG_MLDSA_CTRL                                                                        (32'h10)
`define MLDSA_REG_MLDSA_CTRL_CTRL_LOW                                                               (0)
`define MLDSA_REG_MLDSA_CTRL_CTRL_MASK                                                              (32'h7)
`define MLDSA_REG_MLDSA_CTRL_ZEROIZE_LOW                                                            (3)
`define MLDSA_REG_MLDSA_CTRL_ZEROIZE_MASK                                                           (32'h8)
`define CLP_MLDSA_REG_MLDSA_STATUS                                                                  (32'h10030014)
`define MLDSA_REG_MLDSA_STATUS                                                                      (32'h14)
`define MLDSA_REG_MLDSA_STATUS_READY_LOW                                                            (0)
`define MLDSA_REG_MLDSA_STATUS_READY_MASK                                                           (32'h1)
`define MLDSA_REG_MLDSA_STATUS_VALID_LOW                                                            (1)
`define MLDSA_REG_MLDSA_STATUS_VALID_MASK                                                           (32'h2)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_0                                                               (32'h10030018)
`define MLDSA_REG_MLDSA_ENTROPY_0                                                                   (32'h18)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_1                                                               (32'h1003001c)
`define MLDSA_REG_MLDSA_ENTROPY_1                                                                   (32'h1c)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_2                                                               (32'h10030020)
`define MLDSA_REG_MLDSA_ENTROPY_2                                                                   (32'h20)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_3                                                               (32'h10030024)
`define MLDSA_REG_MLDSA_ENTROPY_3                                                                   (32'h24)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_4                                                               (32'h10030028)
`define MLDSA_REG_MLDSA_ENTROPY_4                                                                   (32'h28)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_5                                                               (32'h1003002c)
`define MLDSA_REG_MLDSA_ENTROPY_5                                                                   (32'h2c)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_6                                                               (32'h10030030)
`define MLDSA_REG_MLDSA_ENTROPY_6                                                                   (32'h30)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_7                                                               (32'h10030034)
`define MLDSA_REG_MLDSA_ENTROPY_7                                                                   (32'h34)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_8                                                               (32'h10030038)
`define MLDSA_REG_MLDSA_ENTROPY_8                                                                   (32'h38)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_9                                                               (32'h1003003c)
`define MLDSA_REG_MLDSA_ENTROPY_9                                                                   (32'h3c)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_10                                                              (32'h10030040)
`define MLDSA_REG_MLDSA_ENTROPY_10                                                                  (32'h40)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_11                                                              (32'h10030044)
`define MLDSA_REG_MLDSA_ENTROPY_11                                                                  (32'h44)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_12                                                              (32'h10030048)
`define MLDSA_REG_MLDSA_ENTROPY_12                                                                  (32'h48)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_13                                                              (32'h1003004c)
`define MLDSA_REG_MLDSA_ENTROPY_13                                                                  (32'h4c)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_14                                                              (32'h10030050)
`define MLDSA_REG_MLDSA_ENTROPY_14                                                                  (32'h50)
`define CLP_MLDSA_REG_MLDSA_ENTROPY_15                                                              (32'h10030054)
`define MLDSA_REG_MLDSA_ENTROPY_15                                                                  (32'h54)
`define CLP_MLDSA_REG_MLDSA_SEED_0                                                                  (32'h10030058)
`define MLDSA_REG_MLDSA_SEED_0                                                                      (32'h58)
`define CLP_MLDSA_REG_MLDSA_SEED_1                                                                  (32'h1003005c)
`define MLDSA_REG_MLDSA_SEED_1                                                                      (32'h5c)
`define CLP_MLDSA_REG_MLDSA_SEED_2                                                                  (32'h10030060)
`define MLDSA_REG_MLDSA_SEED_2                                                                      (32'h60)
`define CLP_MLDSA_REG_MLDSA_SEED_3                                                                  (32'h10030064)
`define MLDSA_REG_MLDSA_SEED_3                                                                      (32'h64)
`define CLP_MLDSA_REG_MLDSA_SEED_4                                                                  (32'h10030068)
`define MLDSA_REG_MLDSA_SEED_4                                                                      (32'h68)
`define CLP_MLDSA_REG_MLDSA_SEED_5                                                                  (32'h1003006c)
`define MLDSA_REG_MLDSA_SEED_5                                                                      (32'h6c)
`define CLP_MLDSA_REG_MLDSA_SEED_6                                                                  (32'h10030070)
`define MLDSA_REG_MLDSA_SEED_6                                                                      (32'h70)
`define CLP_MLDSA_REG_MLDSA_SEED_7                                                                  (32'h10030074)
`define MLDSA_REG_MLDSA_SEED_7                                                                      (32'h74)
`define CLP_MLDSA_REG_MLDSA_SIGN_RND_0                                                              (32'h10030078)
`define MLDSA_REG_MLDSA_SIGN_RND_0                                                                  (32'h78)
`define CLP_MLDSA_REG_MLDSA_SIGN_RND_1                                                              (32'h1003007c)
`define MLDSA_REG_MLDSA_SIGN_RND_1                                                                  (32'h7c)
`define CLP_MLDSA_REG_MLDSA_SIGN_RND_2                                                              (32'h10030080)
`define MLDSA_REG_MLDSA_SIGN_RND_2                                                                  (32'h80)
`define CLP_MLDSA_REG_MLDSA_SIGN_RND_3                                                              (32'h10030084)
`define MLDSA_REG_MLDSA_SIGN_RND_3                                                                  (32'h84)
`define CLP_MLDSA_REG_MLDSA_SIGN_RND_4                                                              (32'h10030088)
`define MLDSA_REG_MLDSA_SIGN_RND_4                                                                  (32'h88)
`define CLP_MLDSA_REG_MLDSA_SIGN_RND_5                                                              (32'h1003008c)
`define MLDSA_REG_MLDSA_SIGN_RND_5                                                                  (32'h8c)
`define CLP_MLDSA_REG_MLDSA_SIGN_RND_6                                                              (32'h10030090)
`define MLDSA_REG_MLDSA_SIGN_RND_6                                                                  (32'h90)
`define CLP_MLDSA_REG_MLDSA_SIGN_RND_7                                                              (32'h10030094)
`define MLDSA_REG_MLDSA_SIGN_RND_7                                                                  (32'h94)
`define CLP_MLDSA_REG_MLDSA_MSG_0                                                                   (32'h10030098)
`define MLDSA_REG_MLDSA_MSG_0                                                                       (32'h98)
`define CLP_MLDSA_REG_MLDSA_MSG_1                                                                   (32'h1003009c)
`define MLDSA_REG_MLDSA_MSG_1                                                                       (32'h9c)
`define CLP_MLDSA_REG_MLDSA_MSG_2                                                                   (32'h100300a0)
`define MLDSA_REG_MLDSA_MSG_2                                                                       (32'ha0)
`define CLP_MLDSA_REG_MLDSA_MSG_3                                                                   (32'h100300a4)
`define MLDSA_REG_MLDSA_MSG_3                                                                       (32'ha4)
`define CLP_MLDSA_REG_MLDSA_MSG_4                                                                   (32'h100300a8)
`define MLDSA_REG_MLDSA_MSG_4                                                                       (32'ha8)
`define CLP_MLDSA_REG_MLDSA_MSG_5                                                                   (32'h100300ac)
`define MLDSA_REG_MLDSA_MSG_5                                                                       (32'hac)
`define CLP_MLDSA_REG_MLDSA_MSG_6                                                                   (32'h100300b0)
`define MLDSA_REG_MLDSA_MSG_6                                                                       (32'hb0)
`define CLP_MLDSA_REG_MLDSA_MSG_7                                                                   (32'h100300b4)
`define MLDSA_REG_MLDSA_MSG_7                                                                       (32'hb4)
`define CLP_MLDSA_REG_MLDSA_MSG_8                                                                   (32'h100300b8)
`define MLDSA_REG_MLDSA_MSG_8                                                                       (32'hb8)
`define CLP_MLDSA_REG_MLDSA_MSG_9                                                                   (32'h100300bc)
`define MLDSA_REG_MLDSA_MSG_9                                                                       (32'hbc)
`define CLP_MLDSA_REG_MLDSA_MSG_10                                                                  (32'h100300c0)
`define MLDSA_REG_MLDSA_MSG_10                                                                      (32'hc0)
`define CLP_MLDSA_REG_MLDSA_MSG_11                                                                  (32'h100300c4)
`define MLDSA_REG_MLDSA_MSG_11                                                                      (32'hc4)
`define CLP_MLDSA_REG_MLDSA_MSG_12                                                                  (32'h100300c8)
`define MLDSA_REG_MLDSA_MSG_12                                                                      (32'hc8)
`define CLP_MLDSA_REG_MLDSA_MSG_13                                                                  (32'h100300cc)
`define MLDSA_REG_MLDSA_MSG_13                                                                      (32'hcc)
`define CLP_MLDSA_REG_MLDSA_MSG_14                                                                  (32'h100300d0)
`define MLDSA_REG_MLDSA_MSG_14                                                                      (32'hd0)
`define CLP_MLDSA_REG_MLDSA_MSG_15                                                                  (32'h100300d4)
`define MLDSA_REG_MLDSA_MSG_15                                                                      (32'hd4)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_0                                                            (32'h100300d8)
`define MLDSA_REG_MLDSA_VERIFY_RES_0                                                                (32'hd8)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_1                                                            (32'h100300dc)
`define MLDSA_REG_MLDSA_VERIFY_RES_1                                                                (32'hdc)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_2                                                            (32'h100300e0)
`define MLDSA_REG_MLDSA_VERIFY_RES_2                                                                (32'he0)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_3                                                            (32'h100300e4)
`define MLDSA_REG_MLDSA_VERIFY_RES_3                                                                (32'he4)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_4                                                            (32'h100300e8)
`define MLDSA_REG_MLDSA_VERIFY_RES_4                                                                (32'he8)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_5                                                            (32'h100300ec)
`define MLDSA_REG_MLDSA_VERIFY_RES_5                                                                (32'hec)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_6                                                            (32'h100300f0)
`define MLDSA_REG_MLDSA_VERIFY_RES_6                                                                (32'hf0)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_7                                                            (32'h100300f4)
`define MLDSA_REG_MLDSA_VERIFY_RES_7                                                                (32'hf4)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_8                                                            (32'h100300f8)
`define MLDSA_REG_MLDSA_VERIFY_RES_8                                                                (32'hf8)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_9                                                            (32'h100300fc)
`define MLDSA_REG_MLDSA_VERIFY_RES_9                                                                (32'hfc)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_10                                                           (32'h10030100)
`define MLDSA_REG_MLDSA_VERIFY_RES_10                                                               (32'h100)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_11                                                           (32'h10030104)
`define MLDSA_REG_MLDSA_VERIFY_RES_11                                                               (32'h104)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_12                                                           (32'h10030108)
`define MLDSA_REG_MLDSA_VERIFY_RES_12                                                               (32'h108)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_13                                                           (32'h1003010c)
`define MLDSA_REG_MLDSA_VERIFY_RES_13                                                               (32'h10c)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_14                                                           (32'h10030110)
`define MLDSA_REG_MLDSA_VERIFY_RES_14                                                               (32'h110)
`define CLP_MLDSA_REG_MLDSA_VERIFY_RES_15                                                           (32'h10030114)
`define MLDSA_REG_MLDSA_VERIFY_RES_15                                                               (32'h114)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_0                                                                (32'h10030118)
`define MLDSA_REG_MLDSA_PUBKEY_0                                                                    (32'h118)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_1                                                                (32'h1003011c)
`define MLDSA_REG_MLDSA_PUBKEY_1                                                                    (32'h11c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_2                                                                (32'h10030120)
`define MLDSA_REG_MLDSA_PUBKEY_2                                                                    (32'h120)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_3                                                                (32'h10030124)
`define MLDSA_REG_MLDSA_PUBKEY_3                                                                    (32'h124)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_4                                                                (32'h10030128)
`define MLDSA_REG_MLDSA_PUBKEY_4                                                                    (32'h128)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_5                                                                (32'h1003012c)
`define MLDSA_REG_MLDSA_PUBKEY_5                                                                    (32'h12c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_6                                                                (32'h10030130)
`define MLDSA_REG_MLDSA_PUBKEY_6                                                                    (32'h130)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_7                                                                (32'h10030134)
`define MLDSA_REG_MLDSA_PUBKEY_7                                                                    (32'h134)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_8                                                                (32'h10030138)
`define MLDSA_REG_MLDSA_PUBKEY_8                                                                    (32'h138)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_9                                                                (32'h1003013c)
`define MLDSA_REG_MLDSA_PUBKEY_9                                                                    (32'h13c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_10                                                               (32'h10030140)
`define MLDSA_REG_MLDSA_PUBKEY_10                                                                   (32'h140)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_11                                                               (32'h10030144)
`define MLDSA_REG_MLDSA_PUBKEY_11                                                                   (32'h144)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_12                                                               (32'h10030148)
`define MLDSA_REG_MLDSA_PUBKEY_12                                                                   (32'h148)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_13                                                               (32'h1003014c)
`define MLDSA_REG_MLDSA_PUBKEY_13                                                                   (32'h14c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_14                                                               (32'h10030150)
`define MLDSA_REG_MLDSA_PUBKEY_14                                                                   (32'h150)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_15                                                               (32'h10030154)
`define MLDSA_REG_MLDSA_PUBKEY_15                                                                   (32'h154)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_16                                                               (32'h10030158)
`define MLDSA_REG_MLDSA_PUBKEY_16                                                                   (32'h158)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_17                                                               (32'h1003015c)
`define MLDSA_REG_MLDSA_PUBKEY_17                                                                   (32'h15c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_18                                                               (32'h10030160)
`define MLDSA_REG_MLDSA_PUBKEY_18                                                                   (32'h160)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_19                                                               (32'h10030164)
`define MLDSA_REG_MLDSA_PUBKEY_19                                                                   (32'h164)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_20                                                               (32'h10030168)
`define MLDSA_REG_MLDSA_PUBKEY_20                                                                   (32'h168)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_21                                                               (32'h1003016c)
`define MLDSA_REG_MLDSA_PUBKEY_21                                                                   (32'h16c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_22                                                               (32'h10030170)
`define MLDSA_REG_MLDSA_PUBKEY_22                                                                   (32'h170)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_23                                                               (32'h10030174)
`define MLDSA_REG_MLDSA_PUBKEY_23                                                                   (32'h174)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_24                                                               (32'h10030178)
`define MLDSA_REG_MLDSA_PUBKEY_24                                                                   (32'h178)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_25                                                               (32'h1003017c)
`define MLDSA_REG_MLDSA_PUBKEY_25                                                                   (32'h17c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_26                                                               (32'h10030180)
`define MLDSA_REG_MLDSA_PUBKEY_26                                                                   (32'h180)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_27                                                               (32'h10030184)
`define MLDSA_REG_MLDSA_PUBKEY_27                                                                   (32'h184)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_28                                                               (32'h10030188)
`define MLDSA_REG_MLDSA_PUBKEY_28                                                                   (32'h188)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_29                                                               (32'h1003018c)
`define MLDSA_REG_MLDSA_PUBKEY_29                                                                   (32'h18c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_30                                                               (32'h10030190)
`define MLDSA_REG_MLDSA_PUBKEY_30                                                                   (32'h190)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_31                                                               (32'h10030194)
`define MLDSA_REG_MLDSA_PUBKEY_31                                                                   (32'h194)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_32                                                               (32'h10030198)
`define MLDSA_REG_MLDSA_PUBKEY_32                                                                   (32'h198)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_33                                                               (32'h1003019c)
`define MLDSA_REG_MLDSA_PUBKEY_33                                                                   (32'h19c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_34                                                               (32'h100301a0)
`define MLDSA_REG_MLDSA_PUBKEY_34                                                                   (32'h1a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_35                                                               (32'h100301a4)
`define MLDSA_REG_MLDSA_PUBKEY_35                                                                   (32'h1a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_36                                                               (32'h100301a8)
`define MLDSA_REG_MLDSA_PUBKEY_36                                                                   (32'h1a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_37                                                               (32'h100301ac)
`define MLDSA_REG_MLDSA_PUBKEY_37                                                                   (32'h1ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_38                                                               (32'h100301b0)
`define MLDSA_REG_MLDSA_PUBKEY_38                                                                   (32'h1b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_39                                                               (32'h100301b4)
`define MLDSA_REG_MLDSA_PUBKEY_39                                                                   (32'h1b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_40                                                               (32'h100301b8)
`define MLDSA_REG_MLDSA_PUBKEY_40                                                                   (32'h1b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_41                                                               (32'h100301bc)
`define MLDSA_REG_MLDSA_PUBKEY_41                                                                   (32'h1bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_42                                                               (32'h100301c0)
`define MLDSA_REG_MLDSA_PUBKEY_42                                                                   (32'h1c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_43                                                               (32'h100301c4)
`define MLDSA_REG_MLDSA_PUBKEY_43                                                                   (32'h1c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_44                                                               (32'h100301c8)
`define MLDSA_REG_MLDSA_PUBKEY_44                                                                   (32'h1c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_45                                                               (32'h100301cc)
`define MLDSA_REG_MLDSA_PUBKEY_45                                                                   (32'h1cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_46                                                               (32'h100301d0)
`define MLDSA_REG_MLDSA_PUBKEY_46                                                                   (32'h1d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_47                                                               (32'h100301d4)
`define MLDSA_REG_MLDSA_PUBKEY_47                                                                   (32'h1d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_48                                                               (32'h100301d8)
`define MLDSA_REG_MLDSA_PUBKEY_48                                                                   (32'h1d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_49                                                               (32'h100301dc)
`define MLDSA_REG_MLDSA_PUBKEY_49                                                                   (32'h1dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_50                                                               (32'h100301e0)
`define MLDSA_REG_MLDSA_PUBKEY_50                                                                   (32'h1e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_51                                                               (32'h100301e4)
`define MLDSA_REG_MLDSA_PUBKEY_51                                                                   (32'h1e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_52                                                               (32'h100301e8)
`define MLDSA_REG_MLDSA_PUBKEY_52                                                                   (32'h1e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_53                                                               (32'h100301ec)
`define MLDSA_REG_MLDSA_PUBKEY_53                                                                   (32'h1ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_54                                                               (32'h100301f0)
`define MLDSA_REG_MLDSA_PUBKEY_54                                                                   (32'h1f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_55                                                               (32'h100301f4)
`define MLDSA_REG_MLDSA_PUBKEY_55                                                                   (32'h1f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_56                                                               (32'h100301f8)
`define MLDSA_REG_MLDSA_PUBKEY_56                                                                   (32'h1f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_57                                                               (32'h100301fc)
`define MLDSA_REG_MLDSA_PUBKEY_57                                                                   (32'h1fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_58                                                               (32'h10030200)
`define MLDSA_REG_MLDSA_PUBKEY_58                                                                   (32'h200)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_59                                                               (32'h10030204)
`define MLDSA_REG_MLDSA_PUBKEY_59                                                                   (32'h204)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_60                                                               (32'h10030208)
`define MLDSA_REG_MLDSA_PUBKEY_60                                                                   (32'h208)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_61                                                               (32'h1003020c)
`define MLDSA_REG_MLDSA_PUBKEY_61                                                                   (32'h20c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_62                                                               (32'h10030210)
`define MLDSA_REG_MLDSA_PUBKEY_62                                                                   (32'h210)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_63                                                               (32'h10030214)
`define MLDSA_REG_MLDSA_PUBKEY_63                                                                   (32'h214)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_64                                                               (32'h10030218)
`define MLDSA_REG_MLDSA_PUBKEY_64                                                                   (32'h218)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_65                                                               (32'h1003021c)
`define MLDSA_REG_MLDSA_PUBKEY_65                                                                   (32'h21c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_66                                                               (32'h10030220)
`define MLDSA_REG_MLDSA_PUBKEY_66                                                                   (32'h220)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_67                                                               (32'h10030224)
`define MLDSA_REG_MLDSA_PUBKEY_67                                                                   (32'h224)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_68                                                               (32'h10030228)
`define MLDSA_REG_MLDSA_PUBKEY_68                                                                   (32'h228)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_69                                                               (32'h1003022c)
`define MLDSA_REG_MLDSA_PUBKEY_69                                                                   (32'h22c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_70                                                               (32'h10030230)
`define MLDSA_REG_MLDSA_PUBKEY_70                                                                   (32'h230)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_71                                                               (32'h10030234)
`define MLDSA_REG_MLDSA_PUBKEY_71                                                                   (32'h234)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_72                                                               (32'h10030238)
`define MLDSA_REG_MLDSA_PUBKEY_72                                                                   (32'h238)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_73                                                               (32'h1003023c)
`define MLDSA_REG_MLDSA_PUBKEY_73                                                                   (32'h23c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_74                                                               (32'h10030240)
`define MLDSA_REG_MLDSA_PUBKEY_74                                                                   (32'h240)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_75                                                               (32'h10030244)
`define MLDSA_REG_MLDSA_PUBKEY_75                                                                   (32'h244)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_76                                                               (32'h10030248)
`define MLDSA_REG_MLDSA_PUBKEY_76                                                                   (32'h248)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_77                                                               (32'h1003024c)
`define MLDSA_REG_MLDSA_PUBKEY_77                                                                   (32'h24c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_78                                                               (32'h10030250)
`define MLDSA_REG_MLDSA_PUBKEY_78                                                                   (32'h250)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_79                                                               (32'h10030254)
`define MLDSA_REG_MLDSA_PUBKEY_79                                                                   (32'h254)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_80                                                               (32'h10030258)
`define MLDSA_REG_MLDSA_PUBKEY_80                                                                   (32'h258)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_81                                                               (32'h1003025c)
`define MLDSA_REG_MLDSA_PUBKEY_81                                                                   (32'h25c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_82                                                               (32'h10030260)
`define MLDSA_REG_MLDSA_PUBKEY_82                                                                   (32'h260)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_83                                                               (32'h10030264)
`define MLDSA_REG_MLDSA_PUBKEY_83                                                                   (32'h264)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_84                                                               (32'h10030268)
`define MLDSA_REG_MLDSA_PUBKEY_84                                                                   (32'h268)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_85                                                               (32'h1003026c)
`define MLDSA_REG_MLDSA_PUBKEY_85                                                                   (32'h26c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_86                                                               (32'h10030270)
`define MLDSA_REG_MLDSA_PUBKEY_86                                                                   (32'h270)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_87                                                               (32'h10030274)
`define MLDSA_REG_MLDSA_PUBKEY_87                                                                   (32'h274)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_88                                                               (32'h10030278)
`define MLDSA_REG_MLDSA_PUBKEY_88                                                                   (32'h278)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_89                                                               (32'h1003027c)
`define MLDSA_REG_MLDSA_PUBKEY_89                                                                   (32'h27c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_90                                                               (32'h10030280)
`define MLDSA_REG_MLDSA_PUBKEY_90                                                                   (32'h280)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_91                                                               (32'h10030284)
`define MLDSA_REG_MLDSA_PUBKEY_91                                                                   (32'h284)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_92                                                               (32'h10030288)
`define MLDSA_REG_MLDSA_PUBKEY_92                                                                   (32'h288)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_93                                                               (32'h1003028c)
`define MLDSA_REG_MLDSA_PUBKEY_93                                                                   (32'h28c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_94                                                               (32'h10030290)
`define MLDSA_REG_MLDSA_PUBKEY_94                                                                   (32'h290)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_95                                                               (32'h10030294)
`define MLDSA_REG_MLDSA_PUBKEY_95                                                                   (32'h294)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_96                                                               (32'h10030298)
`define MLDSA_REG_MLDSA_PUBKEY_96                                                                   (32'h298)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_97                                                               (32'h1003029c)
`define MLDSA_REG_MLDSA_PUBKEY_97                                                                   (32'h29c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_98                                                               (32'h100302a0)
`define MLDSA_REG_MLDSA_PUBKEY_98                                                                   (32'h2a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_99                                                               (32'h100302a4)
`define MLDSA_REG_MLDSA_PUBKEY_99                                                                   (32'h2a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_100                                                              (32'h100302a8)
`define MLDSA_REG_MLDSA_PUBKEY_100                                                                  (32'h2a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_101                                                              (32'h100302ac)
`define MLDSA_REG_MLDSA_PUBKEY_101                                                                  (32'h2ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_102                                                              (32'h100302b0)
`define MLDSA_REG_MLDSA_PUBKEY_102                                                                  (32'h2b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_103                                                              (32'h100302b4)
`define MLDSA_REG_MLDSA_PUBKEY_103                                                                  (32'h2b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_104                                                              (32'h100302b8)
`define MLDSA_REG_MLDSA_PUBKEY_104                                                                  (32'h2b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_105                                                              (32'h100302bc)
`define MLDSA_REG_MLDSA_PUBKEY_105                                                                  (32'h2bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_106                                                              (32'h100302c0)
`define MLDSA_REG_MLDSA_PUBKEY_106                                                                  (32'h2c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_107                                                              (32'h100302c4)
`define MLDSA_REG_MLDSA_PUBKEY_107                                                                  (32'h2c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_108                                                              (32'h100302c8)
`define MLDSA_REG_MLDSA_PUBKEY_108                                                                  (32'h2c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_109                                                              (32'h100302cc)
`define MLDSA_REG_MLDSA_PUBKEY_109                                                                  (32'h2cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_110                                                              (32'h100302d0)
`define MLDSA_REG_MLDSA_PUBKEY_110                                                                  (32'h2d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_111                                                              (32'h100302d4)
`define MLDSA_REG_MLDSA_PUBKEY_111                                                                  (32'h2d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_112                                                              (32'h100302d8)
`define MLDSA_REG_MLDSA_PUBKEY_112                                                                  (32'h2d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_113                                                              (32'h100302dc)
`define MLDSA_REG_MLDSA_PUBKEY_113                                                                  (32'h2dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_114                                                              (32'h100302e0)
`define MLDSA_REG_MLDSA_PUBKEY_114                                                                  (32'h2e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_115                                                              (32'h100302e4)
`define MLDSA_REG_MLDSA_PUBKEY_115                                                                  (32'h2e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_116                                                              (32'h100302e8)
`define MLDSA_REG_MLDSA_PUBKEY_116                                                                  (32'h2e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_117                                                              (32'h100302ec)
`define MLDSA_REG_MLDSA_PUBKEY_117                                                                  (32'h2ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_118                                                              (32'h100302f0)
`define MLDSA_REG_MLDSA_PUBKEY_118                                                                  (32'h2f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_119                                                              (32'h100302f4)
`define MLDSA_REG_MLDSA_PUBKEY_119                                                                  (32'h2f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_120                                                              (32'h100302f8)
`define MLDSA_REG_MLDSA_PUBKEY_120                                                                  (32'h2f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_121                                                              (32'h100302fc)
`define MLDSA_REG_MLDSA_PUBKEY_121                                                                  (32'h2fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_122                                                              (32'h10030300)
`define MLDSA_REG_MLDSA_PUBKEY_122                                                                  (32'h300)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_123                                                              (32'h10030304)
`define MLDSA_REG_MLDSA_PUBKEY_123                                                                  (32'h304)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_124                                                              (32'h10030308)
`define MLDSA_REG_MLDSA_PUBKEY_124                                                                  (32'h308)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_125                                                              (32'h1003030c)
`define MLDSA_REG_MLDSA_PUBKEY_125                                                                  (32'h30c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_126                                                              (32'h10030310)
`define MLDSA_REG_MLDSA_PUBKEY_126                                                                  (32'h310)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_127                                                              (32'h10030314)
`define MLDSA_REG_MLDSA_PUBKEY_127                                                                  (32'h314)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_128                                                              (32'h10030318)
`define MLDSA_REG_MLDSA_PUBKEY_128                                                                  (32'h318)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_129                                                              (32'h1003031c)
`define MLDSA_REG_MLDSA_PUBKEY_129                                                                  (32'h31c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_130                                                              (32'h10030320)
`define MLDSA_REG_MLDSA_PUBKEY_130                                                                  (32'h320)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_131                                                              (32'h10030324)
`define MLDSA_REG_MLDSA_PUBKEY_131                                                                  (32'h324)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_132                                                              (32'h10030328)
`define MLDSA_REG_MLDSA_PUBKEY_132                                                                  (32'h328)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_133                                                              (32'h1003032c)
`define MLDSA_REG_MLDSA_PUBKEY_133                                                                  (32'h32c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_134                                                              (32'h10030330)
`define MLDSA_REG_MLDSA_PUBKEY_134                                                                  (32'h330)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_135                                                              (32'h10030334)
`define MLDSA_REG_MLDSA_PUBKEY_135                                                                  (32'h334)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_136                                                              (32'h10030338)
`define MLDSA_REG_MLDSA_PUBKEY_136                                                                  (32'h338)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_137                                                              (32'h1003033c)
`define MLDSA_REG_MLDSA_PUBKEY_137                                                                  (32'h33c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_138                                                              (32'h10030340)
`define MLDSA_REG_MLDSA_PUBKEY_138                                                                  (32'h340)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_139                                                              (32'h10030344)
`define MLDSA_REG_MLDSA_PUBKEY_139                                                                  (32'h344)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_140                                                              (32'h10030348)
`define MLDSA_REG_MLDSA_PUBKEY_140                                                                  (32'h348)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_141                                                              (32'h1003034c)
`define MLDSA_REG_MLDSA_PUBKEY_141                                                                  (32'h34c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_142                                                              (32'h10030350)
`define MLDSA_REG_MLDSA_PUBKEY_142                                                                  (32'h350)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_143                                                              (32'h10030354)
`define MLDSA_REG_MLDSA_PUBKEY_143                                                                  (32'h354)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_144                                                              (32'h10030358)
`define MLDSA_REG_MLDSA_PUBKEY_144                                                                  (32'h358)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_145                                                              (32'h1003035c)
`define MLDSA_REG_MLDSA_PUBKEY_145                                                                  (32'h35c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_146                                                              (32'h10030360)
`define MLDSA_REG_MLDSA_PUBKEY_146                                                                  (32'h360)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_147                                                              (32'h10030364)
`define MLDSA_REG_MLDSA_PUBKEY_147                                                                  (32'h364)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_148                                                              (32'h10030368)
`define MLDSA_REG_MLDSA_PUBKEY_148                                                                  (32'h368)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_149                                                              (32'h1003036c)
`define MLDSA_REG_MLDSA_PUBKEY_149                                                                  (32'h36c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_150                                                              (32'h10030370)
`define MLDSA_REG_MLDSA_PUBKEY_150                                                                  (32'h370)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_151                                                              (32'h10030374)
`define MLDSA_REG_MLDSA_PUBKEY_151                                                                  (32'h374)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_152                                                              (32'h10030378)
`define MLDSA_REG_MLDSA_PUBKEY_152                                                                  (32'h378)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_153                                                              (32'h1003037c)
`define MLDSA_REG_MLDSA_PUBKEY_153                                                                  (32'h37c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_154                                                              (32'h10030380)
`define MLDSA_REG_MLDSA_PUBKEY_154                                                                  (32'h380)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_155                                                              (32'h10030384)
`define MLDSA_REG_MLDSA_PUBKEY_155                                                                  (32'h384)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_156                                                              (32'h10030388)
`define MLDSA_REG_MLDSA_PUBKEY_156                                                                  (32'h388)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_157                                                              (32'h1003038c)
`define MLDSA_REG_MLDSA_PUBKEY_157                                                                  (32'h38c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_158                                                              (32'h10030390)
`define MLDSA_REG_MLDSA_PUBKEY_158                                                                  (32'h390)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_159                                                              (32'h10030394)
`define MLDSA_REG_MLDSA_PUBKEY_159                                                                  (32'h394)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_160                                                              (32'h10030398)
`define MLDSA_REG_MLDSA_PUBKEY_160                                                                  (32'h398)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_161                                                              (32'h1003039c)
`define MLDSA_REG_MLDSA_PUBKEY_161                                                                  (32'h39c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_162                                                              (32'h100303a0)
`define MLDSA_REG_MLDSA_PUBKEY_162                                                                  (32'h3a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_163                                                              (32'h100303a4)
`define MLDSA_REG_MLDSA_PUBKEY_163                                                                  (32'h3a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_164                                                              (32'h100303a8)
`define MLDSA_REG_MLDSA_PUBKEY_164                                                                  (32'h3a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_165                                                              (32'h100303ac)
`define MLDSA_REG_MLDSA_PUBKEY_165                                                                  (32'h3ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_166                                                              (32'h100303b0)
`define MLDSA_REG_MLDSA_PUBKEY_166                                                                  (32'h3b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_167                                                              (32'h100303b4)
`define MLDSA_REG_MLDSA_PUBKEY_167                                                                  (32'h3b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_168                                                              (32'h100303b8)
`define MLDSA_REG_MLDSA_PUBKEY_168                                                                  (32'h3b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_169                                                              (32'h100303bc)
`define MLDSA_REG_MLDSA_PUBKEY_169                                                                  (32'h3bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_170                                                              (32'h100303c0)
`define MLDSA_REG_MLDSA_PUBKEY_170                                                                  (32'h3c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_171                                                              (32'h100303c4)
`define MLDSA_REG_MLDSA_PUBKEY_171                                                                  (32'h3c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_172                                                              (32'h100303c8)
`define MLDSA_REG_MLDSA_PUBKEY_172                                                                  (32'h3c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_173                                                              (32'h100303cc)
`define MLDSA_REG_MLDSA_PUBKEY_173                                                                  (32'h3cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_174                                                              (32'h100303d0)
`define MLDSA_REG_MLDSA_PUBKEY_174                                                                  (32'h3d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_175                                                              (32'h100303d4)
`define MLDSA_REG_MLDSA_PUBKEY_175                                                                  (32'h3d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_176                                                              (32'h100303d8)
`define MLDSA_REG_MLDSA_PUBKEY_176                                                                  (32'h3d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_177                                                              (32'h100303dc)
`define MLDSA_REG_MLDSA_PUBKEY_177                                                                  (32'h3dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_178                                                              (32'h100303e0)
`define MLDSA_REG_MLDSA_PUBKEY_178                                                                  (32'h3e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_179                                                              (32'h100303e4)
`define MLDSA_REG_MLDSA_PUBKEY_179                                                                  (32'h3e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_180                                                              (32'h100303e8)
`define MLDSA_REG_MLDSA_PUBKEY_180                                                                  (32'h3e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_181                                                              (32'h100303ec)
`define MLDSA_REG_MLDSA_PUBKEY_181                                                                  (32'h3ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_182                                                              (32'h100303f0)
`define MLDSA_REG_MLDSA_PUBKEY_182                                                                  (32'h3f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_183                                                              (32'h100303f4)
`define MLDSA_REG_MLDSA_PUBKEY_183                                                                  (32'h3f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_184                                                              (32'h100303f8)
`define MLDSA_REG_MLDSA_PUBKEY_184                                                                  (32'h3f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_185                                                              (32'h100303fc)
`define MLDSA_REG_MLDSA_PUBKEY_185                                                                  (32'h3fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_186                                                              (32'h10030400)
`define MLDSA_REG_MLDSA_PUBKEY_186                                                                  (32'h400)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_187                                                              (32'h10030404)
`define MLDSA_REG_MLDSA_PUBKEY_187                                                                  (32'h404)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_188                                                              (32'h10030408)
`define MLDSA_REG_MLDSA_PUBKEY_188                                                                  (32'h408)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_189                                                              (32'h1003040c)
`define MLDSA_REG_MLDSA_PUBKEY_189                                                                  (32'h40c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_190                                                              (32'h10030410)
`define MLDSA_REG_MLDSA_PUBKEY_190                                                                  (32'h410)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_191                                                              (32'h10030414)
`define MLDSA_REG_MLDSA_PUBKEY_191                                                                  (32'h414)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_192                                                              (32'h10030418)
`define MLDSA_REG_MLDSA_PUBKEY_192                                                                  (32'h418)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_193                                                              (32'h1003041c)
`define MLDSA_REG_MLDSA_PUBKEY_193                                                                  (32'h41c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_194                                                              (32'h10030420)
`define MLDSA_REG_MLDSA_PUBKEY_194                                                                  (32'h420)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_195                                                              (32'h10030424)
`define MLDSA_REG_MLDSA_PUBKEY_195                                                                  (32'h424)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_196                                                              (32'h10030428)
`define MLDSA_REG_MLDSA_PUBKEY_196                                                                  (32'h428)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_197                                                              (32'h1003042c)
`define MLDSA_REG_MLDSA_PUBKEY_197                                                                  (32'h42c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_198                                                              (32'h10030430)
`define MLDSA_REG_MLDSA_PUBKEY_198                                                                  (32'h430)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_199                                                              (32'h10030434)
`define MLDSA_REG_MLDSA_PUBKEY_199                                                                  (32'h434)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_200                                                              (32'h10030438)
`define MLDSA_REG_MLDSA_PUBKEY_200                                                                  (32'h438)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_201                                                              (32'h1003043c)
`define MLDSA_REG_MLDSA_PUBKEY_201                                                                  (32'h43c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_202                                                              (32'h10030440)
`define MLDSA_REG_MLDSA_PUBKEY_202                                                                  (32'h440)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_203                                                              (32'h10030444)
`define MLDSA_REG_MLDSA_PUBKEY_203                                                                  (32'h444)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_204                                                              (32'h10030448)
`define MLDSA_REG_MLDSA_PUBKEY_204                                                                  (32'h448)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_205                                                              (32'h1003044c)
`define MLDSA_REG_MLDSA_PUBKEY_205                                                                  (32'h44c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_206                                                              (32'h10030450)
`define MLDSA_REG_MLDSA_PUBKEY_206                                                                  (32'h450)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_207                                                              (32'h10030454)
`define MLDSA_REG_MLDSA_PUBKEY_207                                                                  (32'h454)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_208                                                              (32'h10030458)
`define MLDSA_REG_MLDSA_PUBKEY_208                                                                  (32'h458)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_209                                                              (32'h1003045c)
`define MLDSA_REG_MLDSA_PUBKEY_209                                                                  (32'h45c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_210                                                              (32'h10030460)
`define MLDSA_REG_MLDSA_PUBKEY_210                                                                  (32'h460)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_211                                                              (32'h10030464)
`define MLDSA_REG_MLDSA_PUBKEY_211                                                                  (32'h464)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_212                                                              (32'h10030468)
`define MLDSA_REG_MLDSA_PUBKEY_212                                                                  (32'h468)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_213                                                              (32'h1003046c)
`define MLDSA_REG_MLDSA_PUBKEY_213                                                                  (32'h46c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_214                                                              (32'h10030470)
`define MLDSA_REG_MLDSA_PUBKEY_214                                                                  (32'h470)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_215                                                              (32'h10030474)
`define MLDSA_REG_MLDSA_PUBKEY_215                                                                  (32'h474)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_216                                                              (32'h10030478)
`define MLDSA_REG_MLDSA_PUBKEY_216                                                                  (32'h478)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_217                                                              (32'h1003047c)
`define MLDSA_REG_MLDSA_PUBKEY_217                                                                  (32'h47c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_218                                                              (32'h10030480)
`define MLDSA_REG_MLDSA_PUBKEY_218                                                                  (32'h480)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_219                                                              (32'h10030484)
`define MLDSA_REG_MLDSA_PUBKEY_219                                                                  (32'h484)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_220                                                              (32'h10030488)
`define MLDSA_REG_MLDSA_PUBKEY_220                                                                  (32'h488)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_221                                                              (32'h1003048c)
`define MLDSA_REG_MLDSA_PUBKEY_221                                                                  (32'h48c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_222                                                              (32'h10030490)
`define MLDSA_REG_MLDSA_PUBKEY_222                                                                  (32'h490)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_223                                                              (32'h10030494)
`define MLDSA_REG_MLDSA_PUBKEY_223                                                                  (32'h494)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_224                                                              (32'h10030498)
`define MLDSA_REG_MLDSA_PUBKEY_224                                                                  (32'h498)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_225                                                              (32'h1003049c)
`define MLDSA_REG_MLDSA_PUBKEY_225                                                                  (32'h49c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_226                                                              (32'h100304a0)
`define MLDSA_REG_MLDSA_PUBKEY_226                                                                  (32'h4a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_227                                                              (32'h100304a4)
`define MLDSA_REG_MLDSA_PUBKEY_227                                                                  (32'h4a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_228                                                              (32'h100304a8)
`define MLDSA_REG_MLDSA_PUBKEY_228                                                                  (32'h4a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_229                                                              (32'h100304ac)
`define MLDSA_REG_MLDSA_PUBKEY_229                                                                  (32'h4ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_230                                                              (32'h100304b0)
`define MLDSA_REG_MLDSA_PUBKEY_230                                                                  (32'h4b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_231                                                              (32'h100304b4)
`define MLDSA_REG_MLDSA_PUBKEY_231                                                                  (32'h4b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_232                                                              (32'h100304b8)
`define MLDSA_REG_MLDSA_PUBKEY_232                                                                  (32'h4b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_233                                                              (32'h100304bc)
`define MLDSA_REG_MLDSA_PUBKEY_233                                                                  (32'h4bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_234                                                              (32'h100304c0)
`define MLDSA_REG_MLDSA_PUBKEY_234                                                                  (32'h4c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_235                                                              (32'h100304c4)
`define MLDSA_REG_MLDSA_PUBKEY_235                                                                  (32'h4c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_236                                                              (32'h100304c8)
`define MLDSA_REG_MLDSA_PUBKEY_236                                                                  (32'h4c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_237                                                              (32'h100304cc)
`define MLDSA_REG_MLDSA_PUBKEY_237                                                                  (32'h4cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_238                                                              (32'h100304d0)
`define MLDSA_REG_MLDSA_PUBKEY_238                                                                  (32'h4d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_239                                                              (32'h100304d4)
`define MLDSA_REG_MLDSA_PUBKEY_239                                                                  (32'h4d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_240                                                              (32'h100304d8)
`define MLDSA_REG_MLDSA_PUBKEY_240                                                                  (32'h4d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_241                                                              (32'h100304dc)
`define MLDSA_REG_MLDSA_PUBKEY_241                                                                  (32'h4dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_242                                                              (32'h100304e0)
`define MLDSA_REG_MLDSA_PUBKEY_242                                                                  (32'h4e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_243                                                              (32'h100304e4)
`define MLDSA_REG_MLDSA_PUBKEY_243                                                                  (32'h4e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_244                                                              (32'h100304e8)
`define MLDSA_REG_MLDSA_PUBKEY_244                                                                  (32'h4e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_245                                                              (32'h100304ec)
`define MLDSA_REG_MLDSA_PUBKEY_245                                                                  (32'h4ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_246                                                              (32'h100304f0)
`define MLDSA_REG_MLDSA_PUBKEY_246                                                                  (32'h4f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_247                                                              (32'h100304f4)
`define MLDSA_REG_MLDSA_PUBKEY_247                                                                  (32'h4f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_248                                                              (32'h100304f8)
`define MLDSA_REG_MLDSA_PUBKEY_248                                                                  (32'h4f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_249                                                              (32'h100304fc)
`define MLDSA_REG_MLDSA_PUBKEY_249                                                                  (32'h4fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_250                                                              (32'h10030500)
`define MLDSA_REG_MLDSA_PUBKEY_250                                                                  (32'h500)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_251                                                              (32'h10030504)
`define MLDSA_REG_MLDSA_PUBKEY_251                                                                  (32'h504)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_252                                                              (32'h10030508)
`define MLDSA_REG_MLDSA_PUBKEY_252                                                                  (32'h508)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_253                                                              (32'h1003050c)
`define MLDSA_REG_MLDSA_PUBKEY_253                                                                  (32'h50c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_254                                                              (32'h10030510)
`define MLDSA_REG_MLDSA_PUBKEY_254                                                                  (32'h510)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_255                                                              (32'h10030514)
`define MLDSA_REG_MLDSA_PUBKEY_255                                                                  (32'h514)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_256                                                              (32'h10030518)
`define MLDSA_REG_MLDSA_PUBKEY_256                                                                  (32'h518)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_257                                                              (32'h1003051c)
`define MLDSA_REG_MLDSA_PUBKEY_257                                                                  (32'h51c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_258                                                              (32'h10030520)
`define MLDSA_REG_MLDSA_PUBKEY_258                                                                  (32'h520)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_259                                                              (32'h10030524)
`define MLDSA_REG_MLDSA_PUBKEY_259                                                                  (32'h524)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_260                                                              (32'h10030528)
`define MLDSA_REG_MLDSA_PUBKEY_260                                                                  (32'h528)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_261                                                              (32'h1003052c)
`define MLDSA_REG_MLDSA_PUBKEY_261                                                                  (32'h52c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_262                                                              (32'h10030530)
`define MLDSA_REG_MLDSA_PUBKEY_262                                                                  (32'h530)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_263                                                              (32'h10030534)
`define MLDSA_REG_MLDSA_PUBKEY_263                                                                  (32'h534)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_264                                                              (32'h10030538)
`define MLDSA_REG_MLDSA_PUBKEY_264                                                                  (32'h538)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_265                                                              (32'h1003053c)
`define MLDSA_REG_MLDSA_PUBKEY_265                                                                  (32'h53c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_266                                                              (32'h10030540)
`define MLDSA_REG_MLDSA_PUBKEY_266                                                                  (32'h540)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_267                                                              (32'h10030544)
`define MLDSA_REG_MLDSA_PUBKEY_267                                                                  (32'h544)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_268                                                              (32'h10030548)
`define MLDSA_REG_MLDSA_PUBKEY_268                                                                  (32'h548)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_269                                                              (32'h1003054c)
`define MLDSA_REG_MLDSA_PUBKEY_269                                                                  (32'h54c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_270                                                              (32'h10030550)
`define MLDSA_REG_MLDSA_PUBKEY_270                                                                  (32'h550)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_271                                                              (32'h10030554)
`define MLDSA_REG_MLDSA_PUBKEY_271                                                                  (32'h554)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_272                                                              (32'h10030558)
`define MLDSA_REG_MLDSA_PUBKEY_272                                                                  (32'h558)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_273                                                              (32'h1003055c)
`define MLDSA_REG_MLDSA_PUBKEY_273                                                                  (32'h55c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_274                                                              (32'h10030560)
`define MLDSA_REG_MLDSA_PUBKEY_274                                                                  (32'h560)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_275                                                              (32'h10030564)
`define MLDSA_REG_MLDSA_PUBKEY_275                                                                  (32'h564)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_276                                                              (32'h10030568)
`define MLDSA_REG_MLDSA_PUBKEY_276                                                                  (32'h568)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_277                                                              (32'h1003056c)
`define MLDSA_REG_MLDSA_PUBKEY_277                                                                  (32'h56c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_278                                                              (32'h10030570)
`define MLDSA_REG_MLDSA_PUBKEY_278                                                                  (32'h570)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_279                                                              (32'h10030574)
`define MLDSA_REG_MLDSA_PUBKEY_279                                                                  (32'h574)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_280                                                              (32'h10030578)
`define MLDSA_REG_MLDSA_PUBKEY_280                                                                  (32'h578)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_281                                                              (32'h1003057c)
`define MLDSA_REG_MLDSA_PUBKEY_281                                                                  (32'h57c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_282                                                              (32'h10030580)
`define MLDSA_REG_MLDSA_PUBKEY_282                                                                  (32'h580)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_283                                                              (32'h10030584)
`define MLDSA_REG_MLDSA_PUBKEY_283                                                                  (32'h584)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_284                                                              (32'h10030588)
`define MLDSA_REG_MLDSA_PUBKEY_284                                                                  (32'h588)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_285                                                              (32'h1003058c)
`define MLDSA_REG_MLDSA_PUBKEY_285                                                                  (32'h58c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_286                                                              (32'h10030590)
`define MLDSA_REG_MLDSA_PUBKEY_286                                                                  (32'h590)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_287                                                              (32'h10030594)
`define MLDSA_REG_MLDSA_PUBKEY_287                                                                  (32'h594)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_288                                                              (32'h10030598)
`define MLDSA_REG_MLDSA_PUBKEY_288                                                                  (32'h598)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_289                                                              (32'h1003059c)
`define MLDSA_REG_MLDSA_PUBKEY_289                                                                  (32'h59c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_290                                                              (32'h100305a0)
`define MLDSA_REG_MLDSA_PUBKEY_290                                                                  (32'h5a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_291                                                              (32'h100305a4)
`define MLDSA_REG_MLDSA_PUBKEY_291                                                                  (32'h5a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_292                                                              (32'h100305a8)
`define MLDSA_REG_MLDSA_PUBKEY_292                                                                  (32'h5a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_293                                                              (32'h100305ac)
`define MLDSA_REG_MLDSA_PUBKEY_293                                                                  (32'h5ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_294                                                              (32'h100305b0)
`define MLDSA_REG_MLDSA_PUBKEY_294                                                                  (32'h5b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_295                                                              (32'h100305b4)
`define MLDSA_REG_MLDSA_PUBKEY_295                                                                  (32'h5b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_296                                                              (32'h100305b8)
`define MLDSA_REG_MLDSA_PUBKEY_296                                                                  (32'h5b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_297                                                              (32'h100305bc)
`define MLDSA_REG_MLDSA_PUBKEY_297                                                                  (32'h5bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_298                                                              (32'h100305c0)
`define MLDSA_REG_MLDSA_PUBKEY_298                                                                  (32'h5c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_299                                                              (32'h100305c4)
`define MLDSA_REG_MLDSA_PUBKEY_299                                                                  (32'h5c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_300                                                              (32'h100305c8)
`define MLDSA_REG_MLDSA_PUBKEY_300                                                                  (32'h5c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_301                                                              (32'h100305cc)
`define MLDSA_REG_MLDSA_PUBKEY_301                                                                  (32'h5cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_302                                                              (32'h100305d0)
`define MLDSA_REG_MLDSA_PUBKEY_302                                                                  (32'h5d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_303                                                              (32'h100305d4)
`define MLDSA_REG_MLDSA_PUBKEY_303                                                                  (32'h5d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_304                                                              (32'h100305d8)
`define MLDSA_REG_MLDSA_PUBKEY_304                                                                  (32'h5d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_305                                                              (32'h100305dc)
`define MLDSA_REG_MLDSA_PUBKEY_305                                                                  (32'h5dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_306                                                              (32'h100305e0)
`define MLDSA_REG_MLDSA_PUBKEY_306                                                                  (32'h5e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_307                                                              (32'h100305e4)
`define MLDSA_REG_MLDSA_PUBKEY_307                                                                  (32'h5e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_308                                                              (32'h100305e8)
`define MLDSA_REG_MLDSA_PUBKEY_308                                                                  (32'h5e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_309                                                              (32'h100305ec)
`define MLDSA_REG_MLDSA_PUBKEY_309                                                                  (32'h5ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_310                                                              (32'h100305f0)
`define MLDSA_REG_MLDSA_PUBKEY_310                                                                  (32'h5f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_311                                                              (32'h100305f4)
`define MLDSA_REG_MLDSA_PUBKEY_311                                                                  (32'h5f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_312                                                              (32'h100305f8)
`define MLDSA_REG_MLDSA_PUBKEY_312                                                                  (32'h5f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_313                                                              (32'h100305fc)
`define MLDSA_REG_MLDSA_PUBKEY_313                                                                  (32'h5fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_314                                                              (32'h10030600)
`define MLDSA_REG_MLDSA_PUBKEY_314                                                                  (32'h600)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_315                                                              (32'h10030604)
`define MLDSA_REG_MLDSA_PUBKEY_315                                                                  (32'h604)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_316                                                              (32'h10030608)
`define MLDSA_REG_MLDSA_PUBKEY_316                                                                  (32'h608)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_317                                                              (32'h1003060c)
`define MLDSA_REG_MLDSA_PUBKEY_317                                                                  (32'h60c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_318                                                              (32'h10030610)
`define MLDSA_REG_MLDSA_PUBKEY_318                                                                  (32'h610)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_319                                                              (32'h10030614)
`define MLDSA_REG_MLDSA_PUBKEY_319                                                                  (32'h614)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_320                                                              (32'h10030618)
`define MLDSA_REG_MLDSA_PUBKEY_320                                                                  (32'h618)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_321                                                              (32'h1003061c)
`define MLDSA_REG_MLDSA_PUBKEY_321                                                                  (32'h61c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_322                                                              (32'h10030620)
`define MLDSA_REG_MLDSA_PUBKEY_322                                                                  (32'h620)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_323                                                              (32'h10030624)
`define MLDSA_REG_MLDSA_PUBKEY_323                                                                  (32'h624)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_324                                                              (32'h10030628)
`define MLDSA_REG_MLDSA_PUBKEY_324                                                                  (32'h628)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_325                                                              (32'h1003062c)
`define MLDSA_REG_MLDSA_PUBKEY_325                                                                  (32'h62c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_326                                                              (32'h10030630)
`define MLDSA_REG_MLDSA_PUBKEY_326                                                                  (32'h630)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_327                                                              (32'h10030634)
`define MLDSA_REG_MLDSA_PUBKEY_327                                                                  (32'h634)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_328                                                              (32'h10030638)
`define MLDSA_REG_MLDSA_PUBKEY_328                                                                  (32'h638)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_329                                                              (32'h1003063c)
`define MLDSA_REG_MLDSA_PUBKEY_329                                                                  (32'h63c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_330                                                              (32'h10030640)
`define MLDSA_REG_MLDSA_PUBKEY_330                                                                  (32'h640)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_331                                                              (32'h10030644)
`define MLDSA_REG_MLDSA_PUBKEY_331                                                                  (32'h644)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_332                                                              (32'h10030648)
`define MLDSA_REG_MLDSA_PUBKEY_332                                                                  (32'h648)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_333                                                              (32'h1003064c)
`define MLDSA_REG_MLDSA_PUBKEY_333                                                                  (32'h64c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_334                                                              (32'h10030650)
`define MLDSA_REG_MLDSA_PUBKEY_334                                                                  (32'h650)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_335                                                              (32'h10030654)
`define MLDSA_REG_MLDSA_PUBKEY_335                                                                  (32'h654)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_336                                                              (32'h10030658)
`define MLDSA_REG_MLDSA_PUBKEY_336                                                                  (32'h658)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_337                                                              (32'h1003065c)
`define MLDSA_REG_MLDSA_PUBKEY_337                                                                  (32'h65c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_338                                                              (32'h10030660)
`define MLDSA_REG_MLDSA_PUBKEY_338                                                                  (32'h660)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_339                                                              (32'h10030664)
`define MLDSA_REG_MLDSA_PUBKEY_339                                                                  (32'h664)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_340                                                              (32'h10030668)
`define MLDSA_REG_MLDSA_PUBKEY_340                                                                  (32'h668)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_341                                                              (32'h1003066c)
`define MLDSA_REG_MLDSA_PUBKEY_341                                                                  (32'h66c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_342                                                              (32'h10030670)
`define MLDSA_REG_MLDSA_PUBKEY_342                                                                  (32'h670)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_343                                                              (32'h10030674)
`define MLDSA_REG_MLDSA_PUBKEY_343                                                                  (32'h674)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_344                                                              (32'h10030678)
`define MLDSA_REG_MLDSA_PUBKEY_344                                                                  (32'h678)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_345                                                              (32'h1003067c)
`define MLDSA_REG_MLDSA_PUBKEY_345                                                                  (32'h67c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_346                                                              (32'h10030680)
`define MLDSA_REG_MLDSA_PUBKEY_346                                                                  (32'h680)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_347                                                              (32'h10030684)
`define MLDSA_REG_MLDSA_PUBKEY_347                                                                  (32'h684)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_348                                                              (32'h10030688)
`define MLDSA_REG_MLDSA_PUBKEY_348                                                                  (32'h688)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_349                                                              (32'h1003068c)
`define MLDSA_REG_MLDSA_PUBKEY_349                                                                  (32'h68c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_350                                                              (32'h10030690)
`define MLDSA_REG_MLDSA_PUBKEY_350                                                                  (32'h690)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_351                                                              (32'h10030694)
`define MLDSA_REG_MLDSA_PUBKEY_351                                                                  (32'h694)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_352                                                              (32'h10030698)
`define MLDSA_REG_MLDSA_PUBKEY_352                                                                  (32'h698)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_353                                                              (32'h1003069c)
`define MLDSA_REG_MLDSA_PUBKEY_353                                                                  (32'h69c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_354                                                              (32'h100306a0)
`define MLDSA_REG_MLDSA_PUBKEY_354                                                                  (32'h6a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_355                                                              (32'h100306a4)
`define MLDSA_REG_MLDSA_PUBKEY_355                                                                  (32'h6a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_356                                                              (32'h100306a8)
`define MLDSA_REG_MLDSA_PUBKEY_356                                                                  (32'h6a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_357                                                              (32'h100306ac)
`define MLDSA_REG_MLDSA_PUBKEY_357                                                                  (32'h6ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_358                                                              (32'h100306b0)
`define MLDSA_REG_MLDSA_PUBKEY_358                                                                  (32'h6b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_359                                                              (32'h100306b4)
`define MLDSA_REG_MLDSA_PUBKEY_359                                                                  (32'h6b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_360                                                              (32'h100306b8)
`define MLDSA_REG_MLDSA_PUBKEY_360                                                                  (32'h6b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_361                                                              (32'h100306bc)
`define MLDSA_REG_MLDSA_PUBKEY_361                                                                  (32'h6bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_362                                                              (32'h100306c0)
`define MLDSA_REG_MLDSA_PUBKEY_362                                                                  (32'h6c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_363                                                              (32'h100306c4)
`define MLDSA_REG_MLDSA_PUBKEY_363                                                                  (32'h6c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_364                                                              (32'h100306c8)
`define MLDSA_REG_MLDSA_PUBKEY_364                                                                  (32'h6c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_365                                                              (32'h100306cc)
`define MLDSA_REG_MLDSA_PUBKEY_365                                                                  (32'h6cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_366                                                              (32'h100306d0)
`define MLDSA_REG_MLDSA_PUBKEY_366                                                                  (32'h6d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_367                                                              (32'h100306d4)
`define MLDSA_REG_MLDSA_PUBKEY_367                                                                  (32'h6d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_368                                                              (32'h100306d8)
`define MLDSA_REG_MLDSA_PUBKEY_368                                                                  (32'h6d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_369                                                              (32'h100306dc)
`define MLDSA_REG_MLDSA_PUBKEY_369                                                                  (32'h6dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_370                                                              (32'h100306e0)
`define MLDSA_REG_MLDSA_PUBKEY_370                                                                  (32'h6e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_371                                                              (32'h100306e4)
`define MLDSA_REG_MLDSA_PUBKEY_371                                                                  (32'h6e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_372                                                              (32'h100306e8)
`define MLDSA_REG_MLDSA_PUBKEY_372                                                                  (32'h6e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_373                                                              (32'h100306ec)
`define MLDSA_REG_MLDSA_PUBKEY_373                                                                  (32'h6ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_374                                                              (32'h100306f0)
`define MLDSA_REG_MLDSA_PUBKEY_374                                                                  (32'h6f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_375                                                              (32'h100306f4)
`define MLDSA_REG_MLDSA_PUBKEY_375                                                                  (32'h6f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_376                                                              (32'h100306f8)
`define MLDSA_REG_MLDSA_PUBKEY_376                                                                  (32'h6f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_377                                                              (32'h100306fc)
`define MLDSA_REG_MLDSA_PUBKEY_377                                                                  (32'h6fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_378                                                              (32'h10030700)
`define MLDSA_REG_MLDSA_PUBKEY_378                                                                  (32'h700)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_379                                                              (32'h10030704)
`define MLDSA_REG_MLDSA_PUBKEY_379                                                                  (32'h704)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_380                                                              (32'h10030708)
`define MLDSA_REG_MLDSA_PUBKEY_380                                                                  (32'h708)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_381                                                              (32'h1003070c)
`define MLDSA_REG_MLDSA_PUBKEY_381                                                                  (32'h70c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_382                                                              (32'h10030710)
`define MLDSA_REG_MLDSA_PUBKEY_382                                                                  (32'h710)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_383                                                              (32'h10030714)
`define MLDSA_REG_MLDSA_PUBKEY_383                                                                  (32'h714)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_384                                                              (32'h10030718)
`define MLDSA_REG_MLDSA_PUBKEY_384                                                                  (32'h718)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_385                                                              (32'h1003071c)
`define MLDSA_REG_MLDSA_PUBKEY_385                                                                  (32'h71c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_386                                                              (32'h10030720)
`define MLDSA_REG_MLDSA_PUBKEY_386                                                                  (32'h720)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_387                                                              (32'h10030724)
`define MLDSA_REG_MLDSA_PUBKEY_387                                                                  (32'h724)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_388                                                              (32'h10030728)
`define MLDSA_REG_MLDSA_PUBKEY_388                                                                  (32'h728)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_389                                                              (32'h1003072c)
`define MLDSA_REG_MLDSA_PUBKEY_389                                                                  (32'h72c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_390                                                              (32'h10030730)
`define MLDSA_REG_MLDSA_PUBKEY_390                                                                  (32'h730)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_391                                                              (32'h10030734)
`define MLDSA_REG_MLDSA_PUBKEY_391                                                                  (32'h734)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_392                                                              (32'h10030738)
`define MLDSA_REG_MLDSA_PUBKEY_392                                                                  (32'h738)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_393                                                              (32'h1003073c)
`define MLDSA_REG_MLDSA_PUBKEY_393                                                                  (32'h73c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_394                                                              (32'h10030740)
`define MLDSA_REG_MLDSA_PUBKEY_394                                                                  (32'h740)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_395                                                              (32'h10030744)
`define MLDSA_REG_MLDSA_PUBKEY_395                                                                  (32'h744)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_396                                                              (32'h10030748)
`define MLDSA_REG_MLDSA_PUBKEY_396                                                                  (32'h748)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_397                                                              (32'h1003074c)
`define MLDSA_REG_MLDSA_PUBKEY_397                                                                  (32'h74c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_398                                                              (32'h10030750)
`define MLDSA_REG_MLDSA_PUBKEY_398                                                                  (32'h750)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_399                                                              (32'h10030754)
`define MLDSA_REG_MLDSA_PUBKEY_399                                                                  (32'h754)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_400                                                              (32'h10030758)
`define MLDSA_REG_MLDSA_PUBKEY_400                                                                  (32'h758)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_401                                                              (32'h1003075c)
`define MLDSA_REG_MLDSA_PUBKEY_401                                                                  (32'h75c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_402                                                              (32'h10030760)
`define MLDSA_REG_MLDSA_PUBKEY_402                                                                  (32'h760)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_403                                                              (32'h10030764)
`define MLDSA_REG_MLDSA_PUBKEY_403                                                                  (32'h764)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_404                                                              (32'h10030768)
`define MLDSA_REG_MLDSA_PUBKEY_404                                                                  (32'h768)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_405                                                              (32'h1003076c)
`define MLDSA_REG_MLDSA_PUBKEY_405                                                                  (32'h76c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_406                                                              (32'h10030770)
`define MLDSA_REG_MLDSA_PUBKEY_406                                                                  (32'h770)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_407                                                              (32'h10030774)
`define MLDSA_REG_MLDSA_PUBKEY_407                                                                  (32'h774)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_408                                                              (32'h10030778)
`define MLDSA_REG_MLDSA_PUBKEY_408                                                                  (32'h778)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_409                                                              (32'h1003077c)
`define MLDSA_REG_MLDSA_PUBKEY_409                                                                  (32'h77c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_410                                                              (32'h10030780)
`define MLDSA_REG_MLDSA_PUBKEY_410                                                                  (32'h780)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_411                                                              (32'h10030784)
`define MLDSA_REG_MLDSA_PUBKEY_411                                                                  (32'h784)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_412                                                              (32'h10030788)
`define MLDSA_REG_MLDSA_PUBKEY_412                                                                  (32'h788)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_413                                                              (32'h1003078c)
`define MLDSA_REG_MLDSA_PUBKEY_413                                                                  (32'h78c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_414                                                              (32'h10030790)
`define MLDSA_REG_MLDSA_PUBKEY_414                                                                  (32'h790)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_415                                                              (32'h10030794)
`define MLDSA_REG_MLDSA_PUBKEY_415                                                                  (32'h794)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_416                                                              (32'h10030798)
`define MLDSA_REG_MLDSA_PUBKEY_416                                                                  (32'h798)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_417                                                              (32'h1003079c)
`define MLDSA_REG_MLDSA_PUBKEY_417                                                                  (32'h79c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_418                                                              (32'h100307a0)
`define MLDSA_REG_MLDSA_PUBKEY_418                                                                  (32'h7a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_419                                                              (32'h100307a4)
`define MLDSA_REG_MLDSA_PUBKEY_419                                                                  (32'h7a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_420                                                              (32'h100307a8)
`define MLDSA_REG_MLDSA_PUBKEY_420                                                                  (32'h7a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_421                                                              (32'h100307ac)
`define MLDSA_REG_MLDSA_PUBKEY_421                                                                  (32'h7ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_422                                                              (32'h100307b0)
`define MLDSA_REG_MLDSA_PUBKEY_422                                                                  (32'h7b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_423                                                              (32'h100307b4)
`define MLDSA_REG_MLDSA_PUBKEY_423                                                                  (32'h7b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_424                                                              (32'h100307b8)
`define MLDSA_REG_MLDSA_PUBKEY_424                                                                  (32'h7b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_425                                                              (32'h100307bc)
`define MLDSA_REG_MLDSA_PUBKEY_425                                                                  (32'h7bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_426                                                              (32'h100307c0)
`define MLDSA_REG_MLDSA_PUBKEY_426                                                                  (32'h7c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_427                                                              (32'h100307c4)
`define MLDSA_REG_MLDSA_PUBKEY_427                                                                  (32'h7c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_428                                                              (32'h100307c8)
`define MLDSA_REG_MLDSA_PUBKEY_428                                                                  (32'h7c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_429                                                              (32'h100307cc)
`define MLDSA_REG_MLDSA_PUBKEY_429                                                                  (32'h7cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_430                                                              (32'h100307d0)
`define MLDSA_REG_MLDSA_PUBKEY_430                                                                  (32'h7d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_431                                                              (32'h100307d4)
`define MLDSA_REG_MLDSA_PUBKEY_431                                                                  (32'h7d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_432                                                              (32'h100307d8)
`define MLDSA_REG_MLDSA_PUBKEY_432                                                                  (32'h7d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_433                                                              (32'h100307dc)
`define MLDSA_REG_MLDSA_PUBKEY_433                                                                  (32'h7dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_434                                                              (32'h100307e0)
`define MLDSA_REG_MLDSA_PUBKEY_434                                                                  (32'h7e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_435                                                              (32'h100307e4)
`define MLDSA_REG_MLDSA_PUBKEY_435                                                                  (32'h7e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_436                                                              (32'h100307e8)
`define MLDSA_REG_MLDSA_PUBKEY_436                                                                  (32'h7e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_437                                                              (32'h100307ec)
`define MLDSA_REG_MLDSA_PUBKEY_437                                                                  (32'h7ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_438                                                              (32'h100307f0)
`define MLDSA_REG_MLDSA_PUBKEY_438                                                                  (32'h7f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_439                                                              (32'h100307f4)
`define MLDSA_REG_MLDSA_PUBKEY_439                                                                  (32'h7f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_440                                                              (32'h100307f8)
`define MLDSA_REG_MLDSA_PUBKEY_440                                                                  (32'h7f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_441                                                              (32'h100307fc)
`define MLDSA_REG_MLDSA_PUBKEY_441                                                                  (32'h7fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_442                                                              (32'h10030800)
`define MLDSA_REG_MLDSA_PUBKEY_442                                                                  (32'h800)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_443                                                              (32'h10030804)
`define MLDSA_REG_MLDSA_PUBKEY_443                                                                  (32'h804)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_444                                                              (32'h10030808)
`define MLDSA_REG_MLDSA_PUBKEY_444                                                                  (32'h808)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_445                                                              (32'h1003080c)
`define MLDSA_REG_MLDSA_PUBKEY_445                                                                  (32'h80c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_446                                                              (32'h10030810)
`define MLDSA_REG_MLDSA_PUBKEY_446                                                                  (32'h810)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_447                                                              (32'h10030814)
`define MLDSA_REG_MLDSA_PUBKEY_447                                                                  (32'h814)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_448                                                              (32'h10030818)
`define MLDSA_REG_MLDSA_PUBKEY_448                                                                  (32'h818)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_449                                                              (32'h1003081c)
`define MLDSA_REG_MLDSA_PUBKEY_449                                                                  (32'h81c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_450                                                              (32'h10030820)
`define MLDSA_REG_MLDSA_PUBKEY_450                                                                  (32'h820)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_451                                                              (32'h10030824)
`define MLDSA_REG_MLDSA_PUBKEY_451                                                                  (32'h824)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_452                                                              (32'h10030828)
`define MLDSA_REG_MLDSA_PUBKEY_452                                                                  (32'h828)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_453                                                              (32'h1003082c)
`define MLDSA_REG_MLDSA_PUBKEY_453                                                                  (32'h82c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_454                                                              (32'h10030830)
`define MLDSA_REG_MLDSA_PUBKEY_454                                                                  (32'h830)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_455                                                              (32'h10030834)
`define MLDSA_REG_MLDSA_PUBKEY_455                                                                  (32'h834)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_456                                                              (32'h10030838)
`define MLDSA_REG_MLDSA_PUBKEY_456                                                                  (32'h838)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_457                                                              (32'h1003083c)
`define MLDSA_REG_MLDSA_PUBKEY_457                                                                  (32'h83c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_458                                                              (32'h10030840)
`define MLDSA_REG_MLDSA_PUBKEY_458                                                                  (32'h840)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_459                                                              (32'h10030844)
`define MLDSA_REG_MLDSA_PUBKEY_459                                                                  (32'h844)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_460                                                              (32'h10030848)
`define MLDSA_REG_MLDSA_PUBKEY_460                                                                  (32'h848)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_461                                                              (32'h1003084c)
`define MLDSA_REG_MLDSA_PUBKEY_461                                                                  (32'h84c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_462                                                              (32'h10030850)
`define MLDSA_REG_MLDSA_PUBKEY_462                                                                  (32'h850)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_463                                                              (32'h10030854)
`define MLDSA_REG_MLDSA_PUBKEY_463                                                                  (32'h854)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_464                                                              (32'h10030858)
`define MLDSA_REG_MLDSA_PUBKEY_464                                                                  (32'h858)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_465                                                              (32'h1003085c)
`define MLDSA_REG_MLDSA_PUBKEY_465                                                                  (32'h85c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_466                                                              (32'h10030860)
`define MLDSA_REG_MLDSA_PUBKEY_466                                                                  (32'h860)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_467                                                              (32'h10030864)
`define MLDSA_REG_MLDSA_PUBKEY_467                                                                  (32'h864)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_468                                                              (32'h10030868)
`define MLDSA_REG_MLDSA_PUBKEY_468                                                                  (32'h868)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_469                                                              (32'h1003086c)
`define MLDSA_REG_MLDSA_PUBKEY_469                                                                  (32'h86c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_470                                                              (32'h10030870)
`define MLDSA_REG_MLDSA_PUBKEY_470                                                                  (32'h870)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_471                                                              (32'h10030874)
`define MLDSA_REG_MLDSA_PUBKEY_471                                                                  (32'h874)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_472                                                              (32'h10030878)
`define MLDSA_REG_MLDSA_PUBKEY_472                                                                  (32'h878)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_473                                                              (32'h1003087c)
`define MLDSA_REG_MLDSA_PUBKEY_473                                                                  (32'h87c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_474                                                              (32'h10030880)
`define MLDSA_REG_MLDSA_PUBKEY_474                                                                  (32'h880)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_475                                                              (32'h10030884)
`define MLDSA_REG_MLDSA_PUBKEY_475                                                                  (32'h884)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_476                                                              (32'h10030888)
`define MLDSA_REG_MLDSA_PUBKEY_476                                                                  (32'h888)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_477                                                              (32'h1003088c)
`define MLDSA_REG_MLDSA_PUBKEY_477                                                                  (32'h88c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_478                                                              (32'h10030890)
`define MLDSA_REG_MLDSA_PUBKEY_478                                                                  (32'h890)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_479                                                              (32'h10030894)
`define MLDSA_REG_MLDSA_PUBKEY_479                                                                  (32'h894)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_480                                                              (32'h10030898)
`define MLDSA_REG_MLDSA_PUBKEY_480                                                                  (32'h898)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_481                                                              (32'h1003089c)
`define MLDSA_REG_MLDSA_PUBKEY_481                                                                  (32'h89c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_482                                                              (32'h100308a0)
`define MLDSA_REG_MLDSA_PUBKEY_482                                                                  (32'h8a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_483                                                              (32'h100308a4)
`define MLDSA_REG_MLDSA_PUBKEY_483                                                                  (32'h8a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_484                                                              (32'h100308a8)
`define MLDSA_REG_MLDSA_PUBKEY_484                                                                  (32'h8a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_485                                                              (32'h100308ac)
`define MLDSA_REG_MLDSA_PUBKEY_485                                                                  (32'h8ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_486                                                              (32'h100308b0)
`define MLDSA_REG_MLDSA_PUBKEY_486                                                                  (32'h8b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_487                                                              (32'h100308b4)
`define MLDSA_REG_MLDSA_PUBKEY_487                                                                  (32'h8b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_488                                                              (32'h100308b8)
`define MLDSA_REG_MLDSA_PUBKEY_488                                                                  (32'h8b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_489                                                              (32'h100308bc)
`define MLDSA_REG_MLDSA_PUBKEY_489                                                                  (32'h8bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_490                                                              (32'h100308c0)
`define MLDSA_REG_MLDSA_PUBKEY_490                                                                  (32'h8c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_491                                                              (32'h100308c4)
`define MLDSA_REG_MLDSA_PUBKEY_491                                                                  (32'h8c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_492                                                              (32'h100308c8)
`define MLDSA_REG_MLDSA_PUBKEY_492                                                                  (32'h8c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_493                                                              (32'h100308cc)
`define MLDSA_REG_MLDSA_PUBKEY_493                                                                  (32'h8cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_494                                                              (32'h100308d0)
`define MLDSA_REG_MLDSA_PUBKEY_494                                                                  (32'h8d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_495                                                              (32'h100308d4)
`define MLDSA_REG_MLDSA_PUBKEY_495                                                                  (32'h8d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_496                                                              (32'h100308d8)
`define MLDSA_REG_MLDSA_PUBKEY_496                                                                  (32'h8d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_497                                                              (32'h100308dc)
`define MLDSA_REG_MLDSA_PUBKEY_497                                                                  (32'h8dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_498                                                              (32'h100308e0)
`define MLDSA_REG_MLDSA_PUBKEY_498                                                                  (32'h8e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_499                                                              (32'h100308e4)
`define MLDSA_REG_MLDSA_PUBKEY_499                                                                  (32'h8e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_500                                                              (32'h100308e8)
`define MLDSA_REG_MLDSA_PUBKEY_500                                                                  (32'h8e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_501                                                              (32'h100308ec)
`define MLDSA_REG_MLDSA_PUBKEY_501                                                                  (32'h8ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_502                                                              (32'h100308f0)
`define MLDSA_REG_MLDSA_PUBKEY_502                                                                  (32'h8f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_503                                                              (32'h100308f4)
`define MLDSA_REG_MLDSA_PUBKEY_503                                                                  (32'h8f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_504                                                              (32'h100308f8)
`define MLDSA_REG_MLDSA_PUBKEY_504                                                                  (32'h8f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_505                                                              (32'h100308fc)
`define MLDSA_REG_MLDSA_PUBKEY_505                                                                  (32'h8fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_506                                                              (32'h10030900)
`define MLDSA_REG_MLDSA_PUBKEY_506                                                                  (32'h900)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_507                                                              (32'h10030904)
`define MLDSA_REG_MLDSA_PUBKEY_507                                                                  (32'h904)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_508                                                              (32'h10030908)
`define MLDSA_REG_MLDSA_PUBKEY_508                                                                  (32'h908)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_509                                                              (32'h1003090c)
`define MLDSA_REG_MLDSA_PUBKEY_509                                                                  (32'h90c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_510                                                              (32'h10030910)
`define MLDSA_REG_MLDSA_PUBKEY_510                                                                  (32'h910)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_511                                                              (32'h10030914)
`define MLDSA_REG_MLDSA_PUBKEY_511                                                                  (32'h914)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_512                                                              (32'h10030918)
`define MLDSA_REG_MLDSA_PUBKEY_512                                                                  (32'h918)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_513                                                              (32'h1003091c)
`define MLDSA_REG_MLDSA_PUBKEY_513                                                                  (32'h91c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_514                                                              (32'h10030920)
`define MLDSA_REG_MLDSA_PUBKEY_514                                                                  (32'h920)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_515                                                              (32'h10030924)
`define MLDSA_REG_MLDSA_PUBKEY_515                                                                  (32'h924)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_516                                                              (32'h10030928)
`define MLDSA_REG_MLDSA_PUBKEY_516                                                                  (32'h928)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_517                                                              (32'h1003092c)
`define MLDSA_REG_MLDSA_PUBKEY_517                                                                  (32'h92c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_518                                                              (32'h10030930)
`define MLDSA_REG_MLDSA_PUBKEY_518                                                                  (32'h930)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_519                                                              (32'h10030934)
`define MLDSA_REG_MLDSA_PUBKEY_519                                                                  (32'h934)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_520                                                              (32'h10030938)
`define MLDSA_REG_MLDSA_PUBKEY_520                                                                  (32'h938)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_521                                                              (32'h1003093c)
`define MLDSA_REG_MLDSA_PUBKEY_521                                                                  (32'h93c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_522                                                              (32'h10030940)
`define MLDSA_REG_MLDSA_PUBKEY_522                                                                  (32'h940)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_523                                                              (32'h10030944)
`define MLDSA_REG_MLDSA_PUBKEY_523                                                                  (32'h944)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_524                                                              (32'h10030948)
`define MLDSA_REG_MLDSA_PUBKEY_524                                                                  (32'h948)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_525                                                              (32'h1003094c)
`define MLDSA_REG_MLDSA_PUBKEY_525                                                                  (32'h94c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_526                                                              (32'h10030950)
`define MLDSA_REG_MLDSA_PUBKEY_526                                                                  (32'h950)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_527                                                              (32'h10030954)
`define MLDSA_REG_MLDSA_PUBKEY_527                                                                  (32'h954)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_528                                                              (32'h10030958)
`define MLDSA_REG_MLDSA_PUBKEY_528                                                                  (32'h958)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_529                                                              (32'h1003095c)
`define MLDSA_REG_MLDSA_PUBKEY_529                                                                  (32'h95c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_530                                                              (32'h10030960)
`define MLDSA_REG_MLDSA_PUBKEY_530                                                                  (32'h960)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_531                                                              (32'h10030964)
`define MLDSA_REG_MLDSA_PUBKEY_531                                                                  (32'h964)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_532                                                              (32'h10030968)
`define MLDSA_REG_MLDSA_PUBKEY_532                                                                  (32'h968)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_533                                                              (32'h1003096c)
`define MLDSA_REG_MLDSA_PUBKEY_533                                                                  (32'h96c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_534                                                              (32'h10030970)
`define MLDSA_REG_MLDSA_PUBKEY_534                                                                  (32'h970)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_535                                                              (32'h10030974)
`define MLDSA_REG_MLDSA_PUBKEY_535                                                                  (32'h974)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_536                                                              (32'h10030978)
`define MLDSA_REG_MLDSA_PUBKEY_536                                                                  (32'h978)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_537                                                              (32'h1003097c)
`define MLDSA_REG_MLDSA_PUBKEY_537                                                                  (32'h97c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_538                                                              (32'h10030980)
`define MLDSA_REG_MLDSA_PUBKEY_538                                                                  (32'h980)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_539                                                              (32'h10030984)
`define MLDSA_REG_MLDSA_PUBKEY_539                                                                  (32'h984)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_540                                                              (32'h10030988)
`define MLDSA_REG_MLDSA_PUBKEY_540                                                                  (32'h988)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_541                                                              (32'h1003098c)
`define MLDSA_REG_MLDSA_PUBKEY_541                                                                  (32'h98c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_542                                                              (32'h10030990)
`define MLDSA_REG_MLDSA_PUBKEY_542                                                                  (32'h990)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_543                                                              (32'h10030994)
`define MLDSA_REG_MLDSA_PUBKEY_543                                                                  (32'h994)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_544                                                              (32'h10030998)
`define MLDSA_REG_MLDSA_PUBKEY_544                                                                  (32'h998)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_545                                                              (32'h1003099c)
`define MLDSA_REG_MLDSA_PUBKEY_545                                                                  (32'h99c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_546                                                              (32'h100309a0)
`define MLDSA_REG_MLDSA_PUBKEY_546                                                                  (32'h9a0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_547                                                              (32'h100309a4)
`define MLDSA_REG_MLDSA_PUBKEY_547                                                                  (32'h9a4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_548                                                              (32'h100309a8)
`define MLDSA_REG_MLDSA_PUBKEY_548                                                                  (32'h9a8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_549                                                              (32'h100309ac)
`define MLDSA_REG_MLDSA_PUBKEY_549                                                                  (32'h9ac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_550                                                              (32'h100309b0)
`define MLDSA_REG_MLDSA_PUBKEY_550                                                                  (32'h9b0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_551                                                              (32'h100309b4)
`define MLDSA_REG_MLDSA_PUBKEY_551                                                                  (32'h9b4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_552                                                              (32'h100309b8)
`define MLDSA_REG_MLDSA_PUBKEY_552                                                                  (32'h9b8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_553                                                              (32'h100309bc)
`define MLDSA_REG_MLDSA_PUBKEY_553                                                                  (32'h9bc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_554                                                              (32'h100309c0)
`define MLDSA_REG_MLDSA_PUBKEY_554                                                                  (32'h9c0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_555                                                              (32'h100309c4)
`define MLDSA_REG_MLDSA_PUBKEY_555                                                                  (32'h9c4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_556                                                              (32'h100309c8)
`define MLDSA_REG_MLDSA_PUBKEY_556                                                                  (32'h9c8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_557                                                              (32'h100309cc)
`define MLDSA_REG_MLDSA_PUBKEY_557                                                                  (32'h9cc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_558                                                              (32'h100309d0)
`define MLDSA_REG_MLDSA_PUBKEY_558                                                                  (32'h9d0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_559                                                              (32'h100309d4)
`define MLDSA_REG_MLDSA_PUBKEY_559                                                                  (32'h9d4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_560                                                              (32'h100309d8)
`define MLDSA_REG_MLDSA_PUBKEY_560                                                                  (32'h9d8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_561                                                              (32'h100309dc)
`define MLDSA_REG_MLDSA_PUBKEY_561                                                                  (32'h9dc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_562                                                              (32'h100309e0)
`define MLDSA_REG_MLDSA_PUBKEY_562                                                                  (32'h9e0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_563                                                              (32'h100309e4)
`define MLDSA_REG_MLDSA_PUBKEY_563                                                                  (32'h9e4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_564                                                              (32'h100309e8)
`define MLDSA_REG_MLDSA_PUBKEY_564                                                                  (32'h9e8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_565                                                              (32'h100309ec)
`define MLDSA_REG_MLDSA_PUBKEY_565                                                                  (32'h9ec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_566                                                              (32'h100309f0)
`define MLDSA_REG_MLDSA_PUBKEY_566                                                                  (32'h9f0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_567                                                              (32'h100309f4)
`define MLDSA_REG_MLDSA_PUBKEY_567                                                                  (32'h9f4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_568                                                              (32'h100309f8)
`define MLDSA_REG_MLDSA_PUBKEY_568                                                                  (32'h9f8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_569                                                              (32'h100309fc)
`define MLDSA_REG_MLDSA_PUBKEY_569                                                                  (32'h9fc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_570                                                              (32'h10030a00)
`define MLDSA_REG_MLDSA_PUBKEY_570                                                                  (32'ha00)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_571                                                              (32'h10030a04)
`define MLDSA_REG_MLDSA_PUBKEY_571                                                                  (32'ha04)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_572                                                              (32'h10030a08)
`define MLDSA_REG_MLDSA_PUBKEY_572                                                                  (32'ha08)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_573                                                              (32'h10030a0c)
`define MLDSA_REG_MLDSA_PUBKEY_573                                                                  (32'ha0c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_574                                                              (32'h10030a10)
`define MLDSA_REG_MLDSA_PUBKEY_574                                                                  (32'ha10)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_575                                                              (32'h10030a14)
`define MLDSA_REG_MLDSA_PUBKEY_575                                                                  (32'ha14)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_576                                                              (32'h10030a18)
`define MLDSA_REG_MLDSA_PUBKEY_576                                                                  (32'ha18)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_577                                                              (32'h10030a1c)
`define MLDSA_REG_MLDSA_PUBKEY_577                                                                  (32'ha1c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_578                                                              (32'h10030a20)
`define MLDSA_REG_MLDSA_PUBKEY_578                                                                  (32'ha20)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_579                                                              (32'h10030a24)
`define MLDSA_REG_MLDSA_PUBKEY_579                                                                  (32'ha24)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_580                                                              (32'h10030a28)
`define MLDSA_REG_MLDSA_PUBKEY_580                                                                  (32'ha28)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_581                                                              (32'h10030a2c)
`define MLDSA_REG_MLDSA_PUBKEY_581                                                                  (32'ha2c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_582                                                              (32'h10030a30)
`define MLDSA_REG_MLDSA_PUBKEY_582                                                                  (32'ha30)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_583                                                              (32'h10030a34)
`define MLDSA_REG_MLDSA_PUBKEY_583                                                                  (32'ha34)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_584                                                              (32'h10030a38)
`define MLDSA_REG_MLDSA_PUBKEY_584                                                                  (32'ha38)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_585                                                              (32'h10030a3c)
`define MLDSA_REG_MLDSA_PUBKEY_585                                                                  (32'ha3c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_586                                                              (32'h10030a40)
`define MLDSA_REG_MLDSA_PUBKEY_586                                                                  (32'ha40)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_587                                                              (32'h10030a44)
`define MLDSA_REG_MLDSA_PUBKEY_587                                                                  (32'ha44)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_588                                                              (32'h10030a48)
`define MLDSA_REG_MLDSA_PUBKEY_588                                                                  (32'ha48)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_589                                                              (32'h10030a4c)
`define MLDSA_REG_MLDSA_PUBKEY_589                                                                  (32'ha4c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_590                                                              (32'h10030a50)
`define MLDSA_REG_MLDSA_PUBKEY_590                                                                  (32'ha50)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_591                                                              (32'h10030a54)
`define MLDSA_REG_MLDSA_PUBKEY_591                                                                  (32'ha54)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_592                                                              (32'h10030a58)
`define MLDSA_REG_MLDSA_PUBKEY_592                                                                  (32'ha58)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_593                                                              (32'h10030a5c)
`define MLDSA_REG_MLDSA_PUBKEY_593                                                                  (32'ha5c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_594                                                              (32'h10030a60)
`define MLDSA_REG_MLDSA_PUBKEY_594                                                                  (32'ha60)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_595                                                              (32'h10030a64)
`define MLDSA_REG_MLDSA_PUBKEY_595                                                                  (32'ha64)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_596                                                              (32'h10030a68)
`define MLDSA_REG_MLDSA_PUBKEY_596                                                                  (32'ha68)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_597                                                              (32'h10030a6c)
`define MLDSA_REG_MLDSA_PUBKEY_597                                                                  (32'ha6c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_598                                                              (32'h10030a70)
`define MLDSA_REG_MLDSA_PUBKEY_598                                                                  (32'ha70)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_599                                                              (32'h10030a74)
`define MLDSA_REG_MLDSA_PUBKEY_599                                                                  (32'ha74)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_600                                                              (32'h10030a78)
`define MLDSA_REG_MLDSA_PUBKEY_600                                                                  (32'ha78)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_601                                                              (32'h10030a7c)
`define MLDSA_REG_MLDSA_PUBKEY_601                                                                  (32'ha7c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_602                                                              (32'h10030a80)
`define MLDSA_REG_MLDSA_PUBKEY_602                                                                  (32'ha80)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_603                                                              (32'h10030a84)
`define MLDSA_REG_MLDSA_PUBKEY_603                                                                  (32'ha84)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_604                                                              (32'h10030a88)
`define MLDSA_REG_MLDSA_PUBKEY_604                                                                  (32'ha88)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_605                                                              (32'h10030a8c)
`define MLDSA_REG_MLDSA_PUBKEY_605                                                                  (32'ha8c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_606                                                              (32'h10030a90)
`define MLDSA_REG_MLDSA_PUBKEY_606                                                                  (32'ha90)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_607                                                              (32'h10030a94)
`define MLDSA_REG_MLDSA_PUBKEY_607                                                                  (32'ha94)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_608                                                              (32'h10030a98)
`define MLDSA_REG_MLDSA_PUBKEY_608                                                                  (32'ha98)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_609                                                              (32'h10030a9c)
`define MLDSA_REG_MLDSA_PUBKEY_609                                                                  (32'ha9c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_610                                                              (32'h10030aa0)
`define MLDSA_REG_MLDSA_PUBKEY_610                                                                  (32'haa0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_611                                                              (32'h10030aa4)
`define MLDSA_REG_MLDSA_PUBKEY_611                                                                  (32'haa4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_612                                                              (32'h10030aa8)
`define MLDSA_REG_MLDSA_PUBKEY_612                                                                  (32'haa8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_613                                                              (32'h10030aac)
`define MLDSA_REG_MLDSA_PUBKEY_613                                                                  (32'haac)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_614                                                              (32'h10030ab0)
`define MLDSA_REG_MLDSA_PUBKEY_614                                                                  (32'hab0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_615                                                              (32'h10030ab4)
`define MLDSA_REG_MLDSA_PUBKEY_615                                                                  (32'hab4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_616                                                              (32'h10030ab8)
`define MLDSA_REG_MLDSA_PUBKEY_616                                                                  (32'hab8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_617                                                              (32'h10030abc)
`define MLDSA_REG_MLDSA_PUBKEY_617                                                                  (32'habc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_618                                                              (32'h10030ac0)
`define MLDSA_REG_MLDSA_PUBKEY_618                                                                  (32'hac0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_619                                                              (32'h10030ac4)
`define MLDSA_REG_MLDSA_PUBKEY_619                                                                  (32'hac4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_620                                                              (32'h10030ac8)
`define MLDSA_REG_MLDSA_PUBKEY_620                                                                  (32'hac8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_621                                                              (32'h10030acc)
`define MLDSA_REG_MLDSA_PUBKEY_621                                                                  (32'hacc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_622                                                              (32'h10030ad0)
`define MLDSA_REG_MLDSA_PUBKEY_622                                                                  (32'had0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_623                                                              (32'h10030ad4)
`define MLDSA_REG_MLDSA_PUBKEY_623                                                                  (32'had4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_624                                                              (32'h10030ad8)
`define MLDSA_REG_MLDSA_PUBKEY_624                                                                  (32'had8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_625                                                              (32'h10030adc)
`define MLDSA_REG_MLDSA_PUBKEY_625                                                                  (32'hadc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_626                                                              (32'h10030ae0)
`define MLDSA_REG_MLDSA_PUBKEY_626                                                                  (32'hae0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_627                                                              (32'h10030ae4)
`define MLDSA_REG_MLDSA_PUBKEY_627                                                                  (32'hae4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_628                                                              (32'h10030ae8)
`define MLDSA_REG_MLDSA_PUBKEY_628                                                                  (32'hae8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_629                                                              (32'h10030aec)
`define MLDSA_REG_MLDSA_PUBKEY_629                                                                  (32'haec)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_630                                                              (32'h10030af0)
`define MLDSA_REG_MLDSA_PUBKEY_630                                                                  (32'haf0)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_631                                                              (32'h10030af4)
`define MLDSA_REG_MLDSA_PUBKEY_631                                                                  (32'haf4)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_632                                                              (32'h10030af8)
`define MLDSA_REG_MLDSA_PUBKEY_632                                                                  (32'haf8)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_633                                                              (32'h10030afc)
`define MLDSA_REG_MLDSA_PUBKEY_633                                                                  (32'hafc)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_634                                                              (32'h10030b00)
`define MLDSA_REG_MLDSA_PUBKEY_634                                                                  (32'hb00)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_635                                                              (32'h10030b04)
`define MLDSA_REG_MLDSA_PUBKEY_635                                                                  (32'hb04)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_636                                                              (32'h10030b08)
`define MLDSA_REG_MLDSA_PUBKEY_636                                                                  (32'hb08)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_637                                                              (32'h10030b0c)
`define MLDSA_REG_MLDSA_PUBKEY_637                                                                  (32'hb0c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_638                                                              (32'h10030b10)
`define MLDSA_REG_MLDSA_PUBKEY_638                                                                  (32'hb10)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_639                                                              (32'h10030b14)
`define MLDSA_REG_MLDSA_PUBKEY_639                                                                  (32'hb14)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_640                                                              (32'h10030b18)
`define MLDSA_REG_MLDSA_PUBKEY_640                                                                  (32'hb18)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_641                                                              (32'h10030b1c)
`define MLDSA_REG_MLDSA_PUBKEY_641                                                                  (32'hb1c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_642                                                              (32'h10030b20)
`define MLDSA_REG_MLDSA_PUBKEY_642                                                                  (32'hb20)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_643                                                              (32'h10030b24)
`define MLDSA_REG_MLDSA_PUBKEY_643                                                                  (32'hb24)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_644                                                              (32'h10030b28)
`define MLDSA_REG_MLDSA_PUBKEY_644                                                                  (32'hb28)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_645                                                              (32'h10030b2c)
`define MLDSA_REG_MLDSA_PUBKEY_645                                                                  (32'hb2c)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_646                                                              (32'h10030b30)
`define MLDSA_REG_MLDSA_PUBKEY_646                                                                  (32'hb30)
`define CLP_MLDSA_REG_MLDSA_PUBKEY_647                                                              (32'h10030b34)
`define MLDSA_REG_MLDSA_PUBKEY_647                                                                  (32'hb34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_0                                                             (32'h10030b38)
`define MLDSA_REG_MLDSA_SIGNATURE_0                                                                 (32'hb38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1                                                             (32'h10030b3c)
`define MLDSA_REG_MLDSA_SIGNATURE_1                                                                 (32'hb3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_2                                                             (32'h10030b40)
`define MLDSA_REG_MLDSA_SIGNATURE_2                                                                 (32'hb40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_3                                                             (32'h10030b44)
`define MLDSA_REG_MLDSA_SIGNATURE_3                                                                 (32'hb44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_4                                                             (32'h10030b48)
`define MLDSA_REG_MLDSA_SIGNATURE_4                                                                 (32'hb48)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_5                                                             (32'h10030b4c)
`define MLDSA_REG_MLDSA_SIGNATURE_5                                                                 (32'hb4c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_6                                                             (32'h10030b50)
`define MLDSA_REG_MLDSA_SIGNATURE_6                                                                 (32'hb50)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_7                                                             (32'h10030b54)
`define MLDSA_REG_MLDSA_SIGNATURE_7                                                                 (32'hb54)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_8                                                             (32'h10030b58)
`define MLDSA_REG_MLDSA_SIGNATURE_8                                                                 (32'hb58)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_9                                                             (32'h10030b5c)
`define MLDSA_REG_MLDSA_SIGNATURE_9                                                                 (32'hb5c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_10                                                            (32'h10030b60)
`define MLDSA_REG_MLDSA_SIGNATURE_10                                                                (32'hb60)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_11                                                            (32'h10030b64)
`define MLDSA_REG_MLDSA_SIGNATURE_11                                                                (32'hb64)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_12                                                            (32'h10030b68)
`define MLDSA_REG_MLDSA_SIGNATURE_12                                                                (32'hb68)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_13                                                            (32'h10030b6c)
`define MLDSA_REG_MLDSA_SIGNATURE_13                                                                (32'hb6c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_14                                                            (32'h10030b70)
`define MLDSA_REG_MLDSA_SIGNATURE_14                                                                (32'hb70)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_15                                                            (32'h10030b74)
`define MLDSA_REG_MLDSA_SIGNATURE_15                                                                (32'hb74)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_16                                                            (32'h10030b78)
`define MLDSA_REG_MLDSA_SIGNATURE_16                                                                (32'hb78)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_17                                                            (32'h10030b7c)
`define MLDSA_REG_MLDSA_SIGNATURE_17                                                                (32'hb7c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_18                                                            (32'h10030b80)
`define MLDSA_REG_MLDSA_SIGNATURE_18                                                                (32'hb80)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_19                                                            (32'h10030b84)
`define MLDSA_REG_MLDSA_SIGNATURE_19                                                                (32'hb84)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_20                                                            (32'h10030b88)
`define MLDSA_REG_MLDSA_SIGNATURE_20                                                                (32'hb88)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_21                                                            (32'h10030b8c)
`define MLDSA_REG_MLDSA_SIGNATURE_21                                                                (32'hb8c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_22                                                            (32'h10030b90)
`define MLDSA_REG_MLDSA_SIGNATURE_22                                                                (32'hb90)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_23                                                            (32'h10030b94)
`define MLDSA_REG_MLDSA_SIGNATURE_23                                                                (32'hb94)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_24                                                            (32'h10030b98)
`define MLDSA_REG_MLDSA_SIGNATURE_24                                                                (32'hb98)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_25                                                            (32'h10030b9c)
`define MLDSA_REG_MLDSA_SIGNATURE_25                                                                (32'hb9c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_26                                                            (32'h10030ba0)
`define MLDSA_REG_MLDSA_SIGNATURE_26                                                                (32'hba0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_27                                                            (32'h10030ba4)
`define MLDSA_REG_MLDSA_SIGNATURE_27                                                                (32'hba4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_28                                                            (32'h10030ba8)
`define MLDSA_REG_MLDSA_SIGNATURE_28                                                                (32'hba8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_29                                                            (32'h10030bac)
`define MLDSA_REG_MLDSA_SIGNATURE_29                                                                (32'hbac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_30                                                            (32'h10030bb0)
`define MLDSA_REG_MLDSA_SIGNATURE_30                                                                (32'hbb0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_31                                                            (32'h10030bb4)
`define MLDSA_REG_MLDSA_SIGNATURE_31                                                                (32'hbb4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_32                                                            (32'h10030bb8)
`define MLDSA_REG_MLDSA_SIGNATURE_32                                                                (32'hbb8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_33                                                            (32'h10030bbc)
`define MLDSA_REG_MLDSA_SIGNATURE_33                                                                (32'hbbc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_34                                                            (32'h10030bc0)
`define MLDSA_REG_MLDSA_SIGNATURE_34                                                                (32'hbc0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_35                                                            (32'h10030bc4)
`define MLDSA_REG_MLDSA_SIGNATURE_35                                                                (32'hbc4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_36                                                            (32'h10030bc8)
`define MLDSA_REG_MLDSA_SIGNATURE_36                                                                (32'hbc8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_37                                                            (32'h10030bcc)
`define MLDSA_REG_MLDSA_SIGNATURE_37                                                                (32'hbcc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_38                                                            (32'h10030bd0)
`define MLDSA_REG_MLDSA_SIGNATURE_38                                                                (32'hbd0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_39                                                            (32'h10030bd4)
`define MLDSA_REG_MLDSA_SIGNATURE_39                                                                (32'hbd4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_40                                                            (32'h10030bd8)
`define MLDSA_REG_MLDSA_SIGNATURE_40                                                                (32'hbd8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_41                                                            (32'h10030bdc)
`define MLDSA_REG_MLDSA_SIGNATURE_41                                                                (32'hbdc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_42                                                            (32'h10030be0)
`define MLDSA_REG_MLDSA_SIGNATURE_42                                                                (32'hbe0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_43                                                            (32'h10030be4)
`define MLDSA_REG_MLDSA_SIGNATURE_43                                                                (32'hbe4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_44                                                            (32'h10030be8)
`define MLDSA_REG_MLDSA_SIGNATURE_44                                                                (32'hbe8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_45                                                            (32'h10030bec)
`define MLDSA_REG_MLDSA_SIGNATURE_45                                                                (32'hbec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_46                                                            (32'h10030bf0)
`define MLDSA_REG_MLDSA_SIGNATURE_46                                                                (32'hbf0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_47                                                            (32'h10030bf4)
`define MLDSA_REG_MLDSA_SIGNATURE_47                                                                (32'hbf4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_48                                                            (32'h10030bf8)
`define MLDSA_REG_MLDSA_SIGNATURE_48                                                                (32'hbf8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_49                                                            (32'h10030bfc)
`define MLDSA_REG_MLDSA_SIGNATURE_49                                                                (32'hbfc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_50                                                            (32'h10030c00)
`define MLDSA_REG_MLDSA_SIGNATURE_50                                                                (32'hc00)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_51                                                            (32'h10030c04)
`define MLDSA_REG_MLDSA_SIGNATURE_51                                                                (32'hc04)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_52                                                            (32'h10030c08)
`define MLDSA_REG_MLDSA_SIGNATURE_52                                                                (32'hc08)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_53                                                            (32'h10030c0c)
`define MLDSA_REG_MLDSA_SIGNATURE_53                                                                (32'hc0c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_54                                                            (32'h10030c10)
`define MLDSA_REG_MLDSA_SIGNATURE_54                                                                (32'hc10)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_55                                                            (32'h10030c14)
`define MLDSA_REG_MLDSA_SIGNATURE_55                                                                (32'hc14)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_56                                                            (32'h10030c18)
`define MLDSA_REG_MLDSA_SIGNATURE_56                                                                (32'hc18)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_57                                                            (32'h10030c1c)
`define MLDSA_REG_MLDSA_SIGNATURE_57                                                                (32'hc1c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_58                                                            (32'h10030c20)
`define MLDSA_REG_MLDSA_SIGNATURE_58                                                                (32'hc20)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_59                                                            (32'h10030c24)
`define MLDSA_REG_MLDSA_SIGNATURE_59                                                                (32'hc24)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_60                                                            (32'h10030c28)
`define MLDSA_REG_MLDSA_SIGNATURE_60                                                                (32'hc28)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_61                                                            (32'h10030c2c)
`define MLDSA_REG_MLDSA_SIGNATURE_61                                                                (32'hc2c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_62                                                            (32'h10030c30)
`define MLDSA_REG_MLDSA_SIGNATURE_62                                                                (32'hc30)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_63                                                            (32'h10030c34)
`define MLDSA_REG_MLDSA_SIGNATURE_63                                                                (32'hc34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_64                                                            (32'h10030c38)
`define MLDSA_REG_MLDSA_SIGNATURE_64                                                                (32'hc38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_65                                                            (32'h10030c3c)
`define MLDSA_REG_MLDSA_SIGNATURE_65                                                                (32'hc3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_66                                                            (32'h10030c40)
`define MLDSA_REG_MLDSA_SIGNATURE_66                                                                (32'hc40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_67                                                            (32'h10030c44)
`define MLDSA_REG_MLDSA_SIGNATURE_67                                                                (32'hc44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_68                                                            (32'h10030c48)
`define MLDSA_REG_MLDSA_SIGNATURE_68                                                                (32'hc48)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_69                                                            (32'h10030c4c)
`define MLDSA_REG_MLDSA_SIGNATURE_69                                                                (32'hc4c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_70                                                            (32'h10030c50)
`define MLDSA_REG_MLDSA_SIGNATURE_70                                                                (32'hc50)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_71                                                            (32'h10030c54)
`define MLDSA_REG_MLDSA_SIGNATURE_71                                                                (32'hc54)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_72                                                            (32'h10030c58)
`define MLDSA_REG_MLDSA_SIGNATURE_72                                                                (32'hc58)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_73                                                            (32'h10030c5c)
`define MLDSA_REG_MLDSA_SIGNATURE_73                                                                (32'hc5c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_74                                                            (32'h10030c60)
`define MLDSA_REG_MLDSA_SIGNATURE_74                                                                (32'hc60)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_75                                                            (32'h10030c64)
`define MLDSA_REG_MLDSA_SIGNATURE_75                                                                (32'hc64)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_76                                                            (32'h10030c68)
`define MLDSA_REG_MLDSA_SIGNATURE_76                                                                (32'hc68)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_77                                                            (32'h10030c6c)
`define MLDSA_REG_MLDSA_SIGNATURE_77                                                                (32'hc6c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_78                                                            (32'h10030c70)
`define MLDSA_REG_MLDSA_SIGNATURE_78                                                                (32'hc70)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_79                                                            (32'h10030c74)
`define MLDSA_REG_MLDSA_SIGNATURE_79                                                                (32'hc74)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_80                                                            (32'h10030c78)
`define MLDSA_REG_MLDSA_SIGNATURE_80                                                                (32'hc78)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_81                                                            (32'h10030c7c)
`define MLDSA_REG_MLDSA_SIGNATURE_81                                                                (32'hc7c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_82                                                            (32'h10030c80)
`define MLDSA_REG_MLDSA_SIGNATURE_82                                                                (32'hc80)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_83                                                            (32'h10030c84)
`define MLDSA_REG_MLDSA_SIGNATURE_83                                                                (32'hc84)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_84                                                            (32'h10030c88)
`define MLDSA_REG_MLDSA_SIGNATURE_84                                                                (32'hc88)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_85                                                            (32'h10030c8c)
`define MLDSA_REG_MLDSA_SIGNATURE_85                                                                (32'hc8c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_86                                                            (32'h10030c90)
`define MLDSA_REG_MLDSA_SIGNATURE_86                                                                (32'hc90)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_87                                                            (32'h10030c94)
`define MLDSA_REG_MLDSA_SIGNATURE_87                                                                (32'hc94)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_88                                                            (32'h10030c98)
`define MLDSA_REG_MLDSA_SIGNATURE_88                                                                (32'hc98)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_89                                                            (32'h10030c9c)
`define MLDSA_REG_MLDSA_SIGNATURE_89                                                                (32'hc9c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_90                                                            (32'h10030ca0)
`define MLDSA_REG_MLDSA_SIGNATURE_90                                                                (32'hca0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_91                                                            (32'h10030ca4)
`define MLDSA_REG_MLDSA_SIGNATURE_91                                                                (32'hca4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_92                                                            (32'h10030ca8)
`define MLDSA_REG_MLDSA_SIGNATURE_92                                                                (32'hca8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_93                                                            (32'h10030cac)
`define MLDSA_REG_MLDSA_SIGNATURE_93                                                                (32'hcac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_94                                                            (32'h10030cb0)
`define MLDSA_REG_MLDSA_SIGNATURE_94                                                                (32'hcb0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_95                                                            (32'h10030cb4)
`define MLDSA_REG_MLDSA_SIGNATURE_95                                                                (32'hcb4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_96                                                            (32'h10030cb8)
`define MLDSA_REG_MLDSA_SIGNATURE_96                                                                (32'hcb8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_97                                                            (32'h10030cbc)
`define MLDSA_REG_MLDSA_SIGNATURE_97                                                                (32'hcbc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_98                                                            (32'h10030cc0)
`define MLDSA_REG_MLDSA_SIGNATURE_98                                                                (32'hcc0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_99                                                            (32'h10030cc4)
`define MLDSA_REG_MLDSA_SIGNATURE_99                                                                (32'hcc4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_100                                                           (32'h10030cc8)
`define MLDSA_REG_MLDSA_SIGNATURE_100                                                               (32'hcc8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_101                                                           (32'h10030ccc)
`define MLDSA_REG_MLDSA_SIGNATURE_101                                                               (32'hccc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_102                                                           (32'h10030cd0)
`define MLDSA_REG_MLDSA_SIGNATURE_102                                                               (32'hcd0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_103                                                           (32'h10030cd4)
`define MLDSA_REG_MLDSA_SIGNATURE_103                                                               (32'hcd4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_104                                                           (32'h10030cd8)
`define MLDSA_REG_MLDSA_SIGNATURE_104                                                               (32'hcd8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_105                                                           (32'h10030cdc)
`define MLDSA_REG_MLDSA_SIGNATURE_105                                                               (32'hcdc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_106                                                           (32'h10030ce0)
`define MLDSA_REG_MLDSA_SIGNATURE_106                                                               (32'hce0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_107                                                           (32'h10030ce4)
`define MLDSA_REG_MLDSA_SIGNATURE_107                                                               (32'hce4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_108                                                           (32'h10030ce8)
`define MLDSA_REG_MLDSA_SIGNATURE_108                                                               (32'hce8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_109                                                           (32'h10030cec)
`define MLDSA_REG_MLDSA_SIGNATURE_109                                                               (32'hcec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_110                                                           (32'h10030cf0)
`define MLDSA_REG_MLDSA_SIGNATURE_110                                                               (32'hcf0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_111                                                           (32'h10030cf4)
`define MLDSA_REG_MLDSA_SIGNATURE_111                                                               (32'hcf4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_112                                                           (32'h10030cf8)
`define MLDSA_REG_MLDSA_SIGNATURE_112                                                               (32'hcf8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_113                                                           (32'h10030cfc)
`define MLDSA_REG_MLDSA_SIGNATURE_113                                                               (32'hcfc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_114                                                           (32'h10030d00)
`define MLDSA_REG_MLDSA_SIGNATURE_114                                                               (32'hd00)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_115                                                           (32'h10030d04)
`define MLDSA_REG_MLDSA_SIGNATURE_115                                                               (32'hd04)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_116                                                           (32'h10030d08)
`define MLDSA_REG_MLDSA_SIGNATURE_116                                                               (32'hd08)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_117                                                           (32'h10030d0c)
`define MLDSA_REG_MLDSA_SIGNATURE_117                                                               (32'hd0c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_118                                                           (32'h10030d10)
`define MLDSA_REG_MLDSA_SIGNATURE_118                                                               (32'hd10)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_119                                                           (32'h10030d14)
`define MLDSA_REG_MLDSA_SIGNATURE_119                                                               (32'hd14)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_120                                                           (32'h10030d18)
`define MLDSA_REG_MLDSA_SIGNATURE_120                                                               (32'hd18)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_121                                                           (32'h10030d1c)
`define MLDSA_REG_MLDSA_SIGNATURE_121                                                               (32'hd1c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_122                                                           (32'h10030d20)
`define MLDSA_REG_MLDSA_SIGNATURE_122                                                               (32'hd20)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_123                                                           (32'h10030d24)
`define MLDSA_REG_MLDSA_SIGNATURE_123                                                               (32'hd24)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_124                                                           (32'h10030d28)
`define MLDSA_REG_MLDSA_SIGNATURE_124                                                               (32'hd28)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_125                                                           (32'h10030d2c)
`define MLDSA_REG_MLDSA_SIGNATURE_125                                                               (32'hd2c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_126                                                           (32'h10030d30)
`define MLDSA_REG_MLDSA_SIGNATURE_126                                                               (32'hd30)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_127                                                           (32'h10030d34)
`define MLDSA_REG_MLDSA_SIGNATURE_127                                                               (32'hd34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_128                                                           (32'h10030d38)
`define MLDSA_REG_MLDSA_SIGNATURE_128                                                               (32'hd38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_129                                                           (32'h10030d3c)
`define MLDSA_REG_MLDSA_SIGNATURE_129                                                               (32'hd3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_130                                                           (32'h10030d40)
`define MLDSA_REG_MLDSA_SIGNATURE_130                                                               (32'hd40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_131                                                           (32'h10030d44)
`define MLDSA_REG_MLDSA_SIGNATURE_131                                                               (32'hd44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_132                                                           (32'h10030d48)
`define MLDSA_REG_MLDSA_SIGNATURE_132                                                               (32'hd48)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_133                                                           (32'h10030d4c)
`define MLDSA_REG_MLDSA_SIGNATURE_133                                                               (32'hd4c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_134                                                           (32'h10030d50)
`define MLDSA_REG_MLDSA_SIGNATURE_134                                                               (32'hd50)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_135                                                           (32'h10030d54)
`define MLDSA_REG_MLDSA_SIGNATURE_135                                                               (32'hd54)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_136                                                           (32'h10030d58)
`define MLDSA_REG_MLDSA_SIGNATURE_136                                                               (32'hd58)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_137                                                           (32'h10030d5c)
`define MLDSA_REG_MLDSA_SIGNATURE_137                                                               (32'hd5c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_138                                                           (32'h10030d60)
`define MLDSA_REG_MLDSA_SIGNATURE_138                                                               (32'hd60)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_139                                                           (32'h10030d64)
`define MLDSA_REG_MLDSA_SIGNATURE_139                                                               (32'hd64)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_140                                                           (32'h10030d68)
`define MLDSA_REG_MLDSA_SIGNATURE_140                                                               (32'hd68)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_141                                                           (32'h10030d6c)
`define MLDSA_REG_MLDSA_SIGNATURE_141                                                               (32'hd6c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_142                                                           (32'h10030d70)
`define MLDSA_REG_MLDSA_SIGNATURE_142                                                               (32'hd70)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_143                                                           (32'h10030d74)
`define MLDSA_REG_MLDSA_SIGNATURE_143                                                               (32'hd74)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_144                                                           (32'h10030d78)
`define MLDSA_REG_MLDSA_SIGNATURE_144                                                               (32'hd78)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_145                                                           (32'h10030d7c)
`define MLDSA_REG_MLDSA_SIGNATURE_145                                                               (32'hd7c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_146                                                           (32'h10030d80)
`define MLDSA_REG_MLDSA_SIGNATURE_146                                                               (32'hd80)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_147                                                           (32'h10030d84)
`define MLDSA_REG_MLDSA_SIGNATURE_147                                                               (32'hd84)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_148                                                           (32'h10030d88)
`define MLDSA_REG_MLDSA_SIGNATURE_148                                                               (32'hd88)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_149                                                           (32'h10030d8c)
`define MLDSA_REG_MLDSA_SIGNATURE_149                                                               (32'hd8c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_150                                                           (32'h10030d90)
`define MLDSA_REG_MLDSA_SIGNATURE_150                                                               (32'hd90)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_151                                                           (32'h10030d94)
`define MLDSA_REG_MLDSA_SIGNATURE_151                                                               (32'hd94)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_152                                                           (32'h10030d98)
`define MLDSA_REG_MLDSA_SIGNATURE_152                                                               (32'hd98)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_153                                                           (32'h10030d9c)
`define MLDSA_REG_MLDSA_SIGNATURE_153                                                               (32'hd9c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_154                                                           (32'h10030da0)
`define MLDSA_REG_MLDSA_SIGNATURE_154                                                               (32'hda0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_155                                                           (32'h10030da4)
`define MLDSA_REG_MLDSA_SIGNATURE_155                                                               (32'hda4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_156                                                           (32'h10030da8)
`define MLDSA_REG_MLDSA_SIGNATURE_156                                                               (32'hda8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_157                                                           (32'h10030dac)
`define MLDSA_REG_MLDSA_SIGNATURE_157                                                               (32'hdac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_158                                                           (32'h10030db0)
`define MLDSA_REG_MLDSA_SIGNATURE_158                                                               (32'hdb0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_159                                                           (32'h10030db4)
`define MLDSA_REG_MLDSA_SIGNATURE_159                                                               (32'hdb4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_160                                                           (32'h10030db8)
`define MLDSA_REG_MLDSA_SIGNATURE_160                                                               (32'hdb8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_161                                                           (32'h10030dbc)
`define MLDSA_REG_MLDSA_SIGNATURE_161                                                               (32'hdbc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_162                                                           (32'h10030dc0)
`define MLDSA_REG_MLDSA_SIGNATURE_162                                                               (32'hdc0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_163                                                           (32'h10030dc4)
`define MLDSA_REG_MLDSA_SIGNATURE_163                                                               (32'hdc4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_164                                                           (32'h10030dc8)
`define MLDSA_REG_MLDSA_SIGNATURE_164                                                               (32'hdc8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_165                                                           (32'h10030dcc)
`define MLDSA_REG_MLDSA_SIGNATURE_165                                                               (32'hdcc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_166                                                           (32'h10030dd0)
`define MLDSA_REG_MLDSA_SIGNATURE_166                                                               (32'hdd0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_167                                                           (32'h10030dd4)
`define MLDSA_REG_MLDSA_SIGNATURE_167                                                               (32'hdd4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_168                                                           (32'h10030dd8)
`define MLDSA_REG_MLDSA_SIGNATURE_168                                                               (32'hdd8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_169                                                           (32'h10030ddc)
`define MLDSA_REG_MLDSA_SIGNATURE_169                                                               (32'hddc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_170                                                           (32'h10030de0)
`define MLDSA_REG_MLDSA_SIGNATURE_170                                                               (32'hde0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_171                                                           (32'h10030de4)
`define MLDSA_REG_MLDSA_SIGNATURE_171                                                               (32'hde4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_172                                                           (32'h10030de8)
`define MLDSA_REG_MLDSA_SIGNATURE_172                                                               (32'hde8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_173                                                           (32'h10030dec)
`define MLDSA_REG_MLDSA_SIGNATURE_173                                                               (32'hdec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_174                                                           (32'h10030df0)
`define MLDSA_REG_MLDSA_SIGNATURE_174                                                               (32'hdf0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_175                                                           (32'h10030df4)
`define MLDSA_REG_MLDSA_SIGNATURE_175                                                               (32'hdf4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_176                                                           (32'h10030df8)
`define MLDSA_REG_MLDSA_SIGNATURE_176                                                               (32'hdf8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_177                                                           (32'h10030dfc)
`define MLDSA_REG_MLDSA_SIGNATURE_177                                                               (32'hdfc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_178                                                           (32'h10030e00)
`define MLDSA_REG_MLDSA_SIGNATURE_178                                                               (32'he00)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_179                                                           (32'h10030e04)
`define MLDSA_REG_MLDSA_SIGNATURE_179                                                               (32'he04)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_180                                                           (32'h10030e08)
`define MLDSA_REG_MLDSA_SIGNATURE_180                                                               (32'he08)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_181                                                           (32'h10030e0c)
`define MLDSA_REG_MLDSA_SIGNATURE_181                                                               (32'he0c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_182                                                           (32'h10030e10)
`define MLDSA_REG_MLDSA_SIGNATURE_182                                                               (32'he10)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_183                                                           (32'h10030e14)
`define MLDSA_REG_MLDSA_SIGNATURE_183                                                               (32'he14)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_184                                                           (32'h10030e18)
`define MLDSA_REG_MLDSA_SIGNATURE_184                                                               (32'he18)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_185                                                           (32'h10030e1c)
`define MLDSA_REG_MLDSA_SIGNATURE_185                                                               (32'he1c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_186                                                           (32'h10030e20)
`define MLDSA_REG_MLDSA_SIGNATURE_186                                                               (32'he20)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_187                                                           (32'h10030e24)
`define MLDSA_REG_MLDSA_SIGNATURE_187                                                               (32'he24)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_188                                                           (32'h10030e28)
`define MLDSA_REG_MLDSA_SIGNATURE_188                                                               (32'he28)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_189                                                           (32'h10030e2c)
`define MLDSA_REG_MLDSA_SIGNATURE_189                                                               (32'he2c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_190                                                           (32'h10030e30)
`define MLDSA_REG_MLDSA_SIGNATURE_190                                                               (32'he30)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_191                                                           (32'h10030e34)
`define MLDSA_REG_MLDSA_SIGNATURE_191                                                               (32'he34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_192                                                           (32'h10030e38)
`define MLDSA_REG_MLDSA_SIGNATURE_192                                                               (32'he38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_193                                                           (32'h10030e3c)
`define MLDSA_REG_MLDSA_SIGNATURE_193                                                               (32'he3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_194                                                           (32'h10030e40)
`define MLDSA_REG_MLDSA_SIGNATURE_194                                                               (32'he40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_195                                                           (32'h10030e44)
`define MLDSA_REG_MLDSA_SIGNATURE_195                                                               (32'he44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_196                                                           (32'h10030e48)
`define MLDSA_REG_MLDSA_SIGNATURE_196                                                               (32'he48)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_197                                                           (32'h10030e4c)
`define MLDSA_REG_MLDSA_SIGNATURE_197                                                               (32'he4c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_198                                                           (32'h10030e50)
`define MLDSA_REG_MLDSA_SIGNATURE_198                                                               (32'he50)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_199                                                           (32'h10030e54)
`define MLDSA_REG_MLDSA_SIGNATURE_199                                                               (32'he54)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_200                                                           (32'h10030e58)
`define MLDSA_REG_MLDSA_SIGNATURE_200                                                               (32'he58)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_201                                                           (32'h10030e5c)
`define MLDSA_REG_MLDSA_SIGNATURE_201                                                               (32'he5c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_202                                                           (32'h10030e60)
`define MLDSA_REG_MLDSA_SIGNATURE_202                                                               (32'he60)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_203                                                           (32'h10030e64)
`define MLDSA_REG_MLDSA_SIGNATURE_203                                                               (32'he64)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_204                                                           (32'h10030e68)
`define MLDSA_REG_MLDSA_SIGNATURE_204                                                               (32'he68)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_205                                                           (32'h10030e6c)
`define MLDSA_REG_MLDSA_SIGNATURE_205                                                               (32'he6c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_206                                                           (32'h10030e70)
`define MLDSA_REG_MLDSA_SIGNATURE_206                                                               (32'he70)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_207                                                           (32'h10030e74)
`define MLDSA_REG_MLDSA_SIGNATURE_207                                                               (32'he74)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_208                                                           (32'h10030e78)
`define MLDSA_REG_MLDSA_SIGNATURE_208                                                               (32'he78)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_209                                                           (32'h10030e7c)
`define MLDSA_REG_MLDSA_SIGNATURE_209                                                               (32'he7c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_210                                                           (32'h10030e80)
`define MLDSA_REG_MLDSA_SIGNATURE_210                                                               (32'he80)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_211                                                           (32'h10030e84)
`define MLDSA_REG_MLDSA_SIGNATURE_211                                                               (32'he84)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_212                                                           (32'h10030e88)
`define MLDSA_REG_MLDSA_SIGNATURE_212                                                               (32'he88)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_213                                                           (32'h10030e8c)
`define MLDSA_REG_MLDSA_SIGNATURE_213                                                               (32'he8c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_214                                                           (32'h10030e90)
`define MLDSA_REG_MLDSA_SIGNATURE_214                                                               (32'he90)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_215                                                           (32'h10030e94)
`define MLDSA_REG_MLDSA_SIGNATURE_215                                                               (32'he94)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_216                                                           (32'h10030e98)
`define MLDSA_REG_MLDSA_SIGNATURE_216                                                               (32'he98)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_217                                                           (32'h10030e9c)
`define MLDSA_REG_MLDSA_SIGNATURE_217                                                               (32'he9c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_218                                                           (32'h10030ea0)
`define MLDSA_REG_MLDSA_SIGNATURE_218                                                               (32'hea0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_219                                                           (32'h10030ea4)
`define MLDSA_REG_MLDSA_SIGNATURE_219                                                               (32'hea4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_220                                                           (32'h10030ea8)
`define MLDSA_REG_MLDSA_SIGNATURE_220                                                               (32'hea8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_221                                                           (32'h10030eac)
`define MLDSA_REG_MLDSA_SIGNATURE_221                                                               (32'heac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_222                                                           (32'h10030eb0)
`define MLDSA_REG_MLDSA_SIGNATURE_222                                                               (32'heb0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_223                                                           (32'h10030eb4)
`define MLDSA_REG_MLDSA_SIGNATURE_223                                                               (32'heb4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_224                                                           (32'h10030eb8)
`define MLDSA_REG_MLDSA_SIGNATURE_224                                                               (32'heb8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_225                                                           (32'h10030ebc)
`define MLDSA_REG_MLDSA_SIGNATURE_225                                                               (32'hebc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_226                                                           (32'h10030ec0)
`define MLDSA_REG_MLDSA_SIGNATURE_226                                                               (32'hec0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_227                                                           (32'h10030ec4)
`define MLDSA_REG_MLDSA_SIGNATURE_227                                                               (32'hec4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_228                                                           (32'h10030ec8)
`define MLDSA_REG_MLDSA_SIGNATURE_228                                                               (32'hec8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_229                                                           (32'h10030ecc)
`define MLDSA_REG_MLDSA_SIGNATURE_229                                                               (32'hecc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_230                                                           (32'h10030ed0)
`define MLDSA_REG_MLDSA_SIGNATURE_230                                                               (32'hed0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_231                                                           (32'h10030ed4)
`define MLDSA_REG_MLDSA_SIGNATURE_231                                                               (32'hed4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_232                                                           (32'h10030ed8)
`define MLDSA_REG_MLDSA_SIGNATURE_232                                                               (32'hed8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_233                                                           (32'h10030edc)
`define MLDSA_REG_MLDSA_SIGNATURE_233                                                               (32'hedc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_234                                                           (32'h10030ee0)
`define MLDSA_REG_MLDSA_SIGNATURE_234                                                               (32'hee0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_235                                                           (32'h10030ee4)
`define MLDSA_REG_MLDSA_SIGNATURE_235                                                               (32'hee4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_236                                                           (32'h10030ee8)
`define MLDSA_REG_MLDSA_SIGNATURE_236                                                               (32'hee8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_237                                                           (32'h10030eec)
`define MLDSA_REG_MLDSA_SIGNATURE_237                                                               (32'heec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_238                                                           (32'h10030ef0)
`define MLDSA_REG_MLDSA_SIGNATURE_238                                                               (32'hef0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_239                                                           (32'h10030ef4)
`define MLDSA_REG_MLDSA_SIGNATURE_239                                                               (32'hef4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_240                                                           (32'h10030ef8)
`define MLDSA_REG_MLDSA_SIGNATURE_240                                                               (32'hef8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_241                                                           (32'h10030efc)
`define MLDSA_REG_MLDSA_SIGNATURE_241                                                               (32'hefc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_242                                                           (32'h10030f00)
`define MLDSA_REG_MLDSA_SIGNATURE_242                                                               (32'hf00)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_243                                                           (32'h10030f04)
`define MLDSA_REG_MLDSA_SIGNATURE_243                                                               (32'hf04)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_244                                                           (32'h10030f08)
`define MLDSA_REG_MLDSA_SIGNATURE_244                                                               (32'hf08)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_245                                                           (32'h10030f0c)
`define MLDSA_REG_MLDSA_SIGNATURE_245                                                               (32'hf0c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_246                                                           (32'h10030f10)
`define MLDSA_REG_MLDSA_SIGNATURE_246                                                               (32'hf10)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_247                                                           (32'h10030f14)
`define MLDSA_REG_MLDSA_SIGNATURE_247                                                               (32'hf14)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_248                                                           (32'h10030f18)
`define MLDSA_REG_MLDSA_SIGNATURE_248                                                               (32'hf18)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_249                                                           (32'h10030f1c)
`define MLDSA_REG_MLDSA_SIGNATURE_249                                                               (32'hf1c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_250                                                           (32'h10030f20)
`define MLDSA_REG_MLDSA_SIGNATURE_250                                                               (32'hf20)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_251                                                           (32'h10030f24)
`define MLDSA_REG_MLDSA_SIGNATURE_251                                                               (32'hf24)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_252                                                           (32'h10030f28)
`define MLDSA_REG_MLDSA_SIGNATURE_252                                                               (32'hf28)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_253                                                           (32'h10030f2c)
`define MLDSA_REG_MLDSA_SIGNATURE_253                                                               (32'hf2c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_254                                                           (32'h10030f30)
`define MLDSA_REG_MLDSA_SIGNATURE_254                                                               (32'hf30)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_255                                                           (32'h10030f34)
`define MLDSA_REG_MLDSA_SIGNATURE_255                                                               (32'hf34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_256                                                           (32'h10030f38)
`define MLDSA_REG_MLDSA_SIGNATURE_256                                                               (32'hf38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_257                                                           (32'h10030f3c)
`define MLDSA_REG_MLDSA_SIGNATURE_257                                                               (32'hf3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_258                                                           (32'h10030f40)
`define MLDSA_REG_MLDSA_SIGNATURE_258                                                               (32'hf40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_259                                                           (32'h10030f44)
`define MLDSA_REG_MLDSA_SIGNATURE_259                                                               (32'hf44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_260                                                           (32'h10030f48)
`define MLDSA_REG_MLDSA_SIGNATURE_260                                                               (32'hf48)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_261                                                           (32'h10030f4c)
`define MLDSA_REG_MLDSA_SIGNATURE_261                                                               (32'hf4c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_262                                                           (32'h10030f50)
`define MLDSA_REG_MLDSA_SIGNATURE_262                                                               (32'hf50)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_263                                                           (32'h10030f54)
`define MLDSA_REG_MLDSA_SIGNATURE_263                                                               (32'hf54)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_264                                                           (32'h10030f58)
`define MLDSA_REG_MLDSA_SIGNATURE_264                                                               (32'hf58)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_265                                                           (32'h10030f5c)
`define MLDSA_REG_MLDSA_SIGNATURE_265                                                               (32'hf5c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_266                                                           (32'h10030f60)
`define MLDSA_REG_MLDSA_SIGNATURE_266                                                               (32'hf60)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_267                                                           (32'h10030f64)
`define MLDSA_REG_MLDSA_SIGNATURE_267                                                               (32'hf64)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_268                                                           (32'h10030f68)
`define MLDSA_REG_MLDSA_SIGNATURE_268                                                               (32'hf68)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_269                                                           (32'h10030f6c)
`define MLDSA_REG_MLDSA_SIGNATURE_269                                                               (32'hf6c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_270                                                           (32'h10030f70)
`define MLDSA_REG_MLDSA_SIGNATURE_270                                                               (32'hf70)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_271                                                           (32'h10030f74)
`define MLDSA_REG_MLDSA_SIGNATURE_271                                                               (32'hf74)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_272                                                           (32'h10030f78)
`define MLDSA_REG_MLDSA_SIGNATURE_272                                                               (32'hf78)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_273                                                           (32'h10030f7c)
`define MLDSA_REG_MLDSA_SIGNATURE_273                                                               (32'hf7c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_274                                                           (32'h10030f80)
`define MLDSA_REG_MLDSA_SIGNATURE_274                                                               (32'hf80)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_275                                                           (32'h10030f84)
`define MLDSA_REG_MLDSA_SIGNATURE_275                                                               (32'hf84)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_276                                                           (32'h10030f88)
`define MLDSA_REG_MLDSA_SIGNATURE_276                                                               (32'hf88)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_277                                                           (32'h10030f8c)
`define MLDSA_REG_MLDSA_SIGNATURE_277                                                               (32'hf8c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_278                                                           (32'h10030f90)
`define MLDSA_REG_MLDSA_SIGNATURE_278                                                               (32'hf90)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_279                                                           (32'h10030f94)
`define MLDSA_REG_MLDSA_SIGNATURE_279                                                               (32'hf94)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_280                                                           (32'h10030f98)
`define MLDSA_REG_MLDSA_SIGNATURE_280                                                               (32'hf98)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_281                                                           (32'h10030f9c)
`define MLDSA_REG_MLDSA_SIGNATURE_281                                                               (32'hf9c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_282                                                           (32'h10030fa0)
`define MLDSA_REG_MLDSA_SIGNATURE_282                                                               (32'hfa0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_283                                                           (32'h10030fa4)
`define MLDSA_REG_MLDSA_SIGNATURE_283                                                               (32'hfa4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_284                                                           (32'h10030fa8)
`define MLDSA_REG_MLDSA_SIGNATURE_284                                                               (32'hfa8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_285                                                           (32'h10030fac)
`define MLDSA_REG_MLDSA_SIGNATURE_285                                                               (32'hfac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_286                                                           (32'h10030fb0)
`define MLDSA_REG_MLDSA_SIGNATURE_286                                                               (32'hfb0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_287                                                           (32'h10030fb4)
`define MLDSA_REG_MLDSA_SIGNATURE_287                                                               (32'hfb4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_288                                                           (32'h10030fb8)
`define MLDSA_REG_MLDSA_SIGNATURE_288                                                               (32'hfb8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_289                                                           (32'h10030fbc)
`define MLDSA_REG_MLDSA_SIGNATURE_289                                                               (32'hfbc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_290                                                           (32'h10030fc0)
`define MLDSA_REG_MLDSA_SIGNATURE_290                                                               (32'hfc0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_291                                                           (32'h10030fc4)
`define MLDSA_REG_MLDSA_SIGNATURE_291                                                               (32'hfc4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_292                                                           (32'h10030fc8)
`define MLDSA_REG_MLDSA_SIGNATURE_292                                                               (32'hfc8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_293                                                           (32'h10030fcc)
`define MLDSA_REG_MLDSA_SIGNATURE_293                                                               (32'hfcc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_294                                                           (32'h10030fd0)
`define MLDSA_REG_MLDSA_SIGNATURE_294                                                               (32'hfd0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_295                                                           (32'h10030fd4)
`define MLDSA_REG_MLDSA_SIGNATURE_295                                                               (32'hfd4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_296                                                           (32'h10030fd8)
`define MLDSA_REG_MLDSA_SIGNATURE_296                                                               (32'hfd8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_297                                                           (32'h10030fdc)
`define MLDSA_REG_MLDSA_SIGNATURE_297                                                               (32'hfdc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_298                                                           (32'h10030fe0)
`define MLDSA_REG_MLDSA_SIGNATURE_298                                                               (32'hfe0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_299                                                           (32'h10030fe4)
`define MLDSA_REG_MLDSA_SIGNATURE_299                                                               (32'hfe4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_300                                                           (32'h10030fe8)
`define MLDSA_REG_MLDSA_SIGNATURE_300                                                               (32'hfe8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_301                                                           (32'h10030fec)
`define MLDSA_REG_MLDSA_SIGNATURE_301                                                               (32'hfec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_302                                                           (32'h10030ff0)
`define MLDSA_REG_MLDSA_SIGNATURE_302                                                               (32'hff0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_303                                                           (32'h10030ff4)
`define MLDSA_REG_MLDSA_SIGNATURE_303                                                               (32'hff4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_304                                                           (32'h10030ff8)
`define MLDSA_REG_MLDSA_SIGNATURE_304                                                               (32'hff8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_305                                                           (32'h10030ffc)
`define MLDSA_REG_MLDSA_SIGNATURE_305                                                               (32'hffc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_306                                                           (32'h10031000)
`define MLDSA_REG_MLDSA_SIGNATURE_306                                                               (32'h1000)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_307                                                           (32'h10031004)
`define MLDSA_REG_MLDSA_SIGNATURE_307                                                               (32'h1004)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_308                                                           (32'h10031008)
`define MLDSA_REG_MLDSA_SIGNATURE_308                                                               (32'h1008)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_309                                                           (32'h1003100c)
`define MLDSA_REG_MLDSA_SIGNATURE_309                                                               (32'h100c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_310                                                           (32'h10031010)
`define MLDSA_REG_MLDSA_SIGNATURE_310                                                               (32'h1010)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_311                                                           (32'h10031014)
`define MLDSA_REG_MLDSA_SIGNATURE_311                                                               (32'h1014)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_312                                                           (32'h10031018)
`define MLDSA_REG_MLDSA_SIGNATURE_312                                                               (32'h1018)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_313                                                           (32'h1003101c)
`define MLDSA_REG_MLDSA_SIGNATURE_313                                                               (32'h101c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_314                                                           (32'h10031020)
`define MLDSA_REG_MLDSA_SIGNATURE_314                                                               (32'h1020)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_315                                                           (32'h10031024)
`define MLDSA_REG_MLDSA_SIGNATURE_315                                                               (32'h1024)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_316                                                           (32'h10031028)
`define MLDSA_REG_MLDSA_SIGNATURE_316                                                               (32'h1028)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_317                                                           (32'h1003102c)
`define MLDSA_REG_MLDSA_SIGNATURE_317                                                               (32'h102c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_318                                                           (32'h10031030)
`define MLDSA_REG_MLDSA_SIGNATURE_318                                                               (32'h1030)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_319                                                           (32'h10031034)
`define MLDSA_REG_MLDSA_SIGNATURE_319                                                               (32'h1034)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_320                                                           (32'h10031038)
`define MLDSA_REG_MLDSA_SIGNATURE_320                                                               (32'h1038)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_321                                                           (32'h1003103c)
`define MLDSA_REG_MLDSA_SIGNATURE_321                                                               (32'h103c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_322                                                           (32'h10031040)
`define MLDSA_REG_MLDSA_SIGNATURE_322                                                               (32'h1040)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_323                                                           (32'h10031044)
`define MLDSA_REG_MLDSA_SIGNATURE_323                                                               (32'h1044)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_324                                                           (32'h10031048)
`define MLDSA_REG_MLDSA_SIGNATURE_324                                                               (32'h1048)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_325                                                           (32'h1003104c)
`define MLDSA_REG_MLDSA_SIGNATURE_325                                                               (32'h104c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_326                                                           (32'h10031050)
`define MLDSA_REG_MLDSA_SIGNATURE_326                                                               (32'h1050)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_327                                                           (32'h10031054)
`define MLDSA_REG_MLDSA_SIGNATURE_327                                                               (32'h1054)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_328                                                           (32'h10031058)
`define MLDSA_REG_MLDSA_SIGNATURE_328                                                               (32'h1058)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_329                                                           (32'h1003105c)
`define MLDSA_REG_MLDSA_SIGNATURE_329                                                               (32'h105c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_330                                                           (32'h10031060)
`define MLDSA_REG_MLDSA_SIGNATURE_330                                                               (32'h1060)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_331                                                           (32'h10031064)
`define MLDSA_REG_MLDSA_SIGNATURE_331                                                               (32'h1064)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_332                                                           (32'h10031068)
`define MLDSA_REG_MLDSA_SIGNATURE_332                                                               (32'h1068)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_333                                                           (32'h1003106c)
`define MLDSA_REG_MLDSA_SIGNATURE_333                                                               (32'h106c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_334                                                           (32'h10031070)
`define MLDSA_REG_MLDSA_SIGNATURE_334                                                               (32'h1070)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_335                                                           (32'h10031074)
`define MLDSA_REG_MLDSA_SIGNATURE_335                                                               (32'h1074)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_336                                                           (32'h10031078)
`define MLDSA_REG_MLDSA_SIGNATURE_336                                                               (32'h1078)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_337                                                           (32'h1003107c)
`define MLDSA_REG_MLDSA_SIGNATURE_337                                                               (32'h107c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_338                                                           (32'h10031080)
`define MLDSA_REG_MLDSA_SIGNATURE_338                                                               (32'h1080)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_339                                                           (32'h10031084)
`define MLDSA_REG_MLDSA_SIGNATURE_339                                                               (32'h1084)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_340                                                           (32'h10031088)
`define MLDSA_REG_MLDSA_SIGNATURE_340                                                               (32'h1088)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_341                                                           (32'h1003108c)
`define MLDSA_REG_MLDSA_SIGNATURE_341                                                               (32'h108c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_342                                                           (32'h10031090)
`define MLDSA_REG_MLDSA_SIGNATURE_342                                                               (32'h1090)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_343                                                           (32'h10031094)
`define MLDSA_REG_MLDSA_SIGNATURE_343                                                               (32'h1094)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_344                                                           (32'h10031098)
`define MLDSA_REG_MLDSA_SIGNATURE_344                                                               (32'h1098)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_345                                                           (32'h1003109c)
`define MLDSA_REG_MLDSA_SIGNATURE_345                                                               (32'h109c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_346                                                           (32'h100310a0)
`define MLDSA_REG_MLDSA_SIGNATURE_346                                                               (32'h10a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_347                                                           (32'h100310a4)
`define MLDSA_REG_MLDSA_SIGNATURE_347                                                               (32'h10a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_348                                                           (32'h100310a8)
`define MLDSA_REG_MLDSA_SIGNATURE_348                                                               (32'h10a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_349                                                           (32'h100310ac)
`define MLDSA_REG_MLDSA_SIGNATURE_349                                                               (32'h10ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_350                                                           (32'h100310b0)
`define MLDSA_REG_MLDSA_SIGNATURE_350                                                               (32'h10b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_351                                                           (32'h100310b4)
`define MLDSA_REG_MLDSA_SIGNATURE_351                                                               (32'h10b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_352                                                           (32'h100310b8)
`define MLDSA_REG_MLDSA_SIGNATURE_352                                                               (32'h10b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_353                                                           (32'h100310bc)
`define MLDSA_REG_MLDSA_SIGNATURE_353                                                               (32'h10bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_354                                                           (32'h100310c0)
`define MLDSA_REG_MLDSA_SIGNATURE_354                                                               (32'h10c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_355                                                           (32'h100310c4)
`define MLDSA_REG_MLDSA_SIGNATURE_355                                                               (32'h10c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_356                                                           (32'h100310c8)
`define MLDSA_REG_MLDSA_SIGNATURE_356                                                               (32'h10c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_357                                                           (32'h100310cc)
`define MLDSA_REG_MLDSA_SIGNATURE_357                                                               (32'h10cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_358                                                           (32'h100310d0)
`define MLDSA_REG_MLDSA_SIGNATURE_358                                                               (32'h10d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_359                                                           (32'h100310d4)
`define MLDSA_REG_MLDSA_SIGNATURE_359                                                               (32'h10d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_360                                                           (32'h100310d8)
`define MLDSA_REG_MLDSA_SIGNATURE_360                                                               (32'h10d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_361                                                           (32'h100310dc)
`define MLDSA_REG_MLDSA_SIGNATURE_361                                                               (32'h10dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_362                                                           (32'h100310e0)
`define MLDSA_REG_MLDSA_SIGNATURE_362                                                               (32'h10e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_363                                                           (32'h100310e4)
`define MLDSA_REG_MLDSA_SIGNATURE_363                                                               (32'h10e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_364                                                           (32'h100310e8)
`define MLDSA_REG_MLDSA_SIGNATURE_364                                                               (32'h10e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_365                                                           (32'h100310ec)
`define MLDSA_REG_MLDSA_SIGNATURE_365                                                               (32'h10ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_366                                                           (32'h100310f0)
`define MLDSA_REG_MLDSA_SIGNATURE_366                                                               (32'h10f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_367                                                           (32'h100310f4)
`define MLDSA_REG_MLDSA_SIGNATURE_367                                                               (32'h10f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_368                                                           (32'h100310f8)
`define MLDSA_REG_MLDSA_SIGNATURE_368                                                               (32'h10f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_369                                                           (32'h100310fc)
`define MLDSA_REG_MLDSA_SIGNATURE_369                                                               (32'h10fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_370                                                           (32'h10031100)
`define MLDSA_REG_MLDSA_SIGNATURE_370                                                               (32'h1100)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_371                                                           (32'h10031104)
`define MLDSA_REG_MLDSA_SIGNATURE_371                                                               (32'h1104)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_372                                                           (32'h10031108)
`define MLDSA_REG_MLDSA_SIGNATURE_372                                                               (32'h1108)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_373                                                           (32'h1003110c)
`define MLDSA_REG_MLDSA_SIGNATURE_373                                                               (32'h110c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_374                                                           (32'h10031110)
`define MLDSA_REG_MLDSA_SIGNATURE_374                                                               (32'h1110)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_375                                                           (32'h10031114)
`define MLDSA_REG_MLDSA_SIGNATURE_375                                                               (32'h1114)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_376                                                           (32'h10031118)
`define MLDSA_REG_MLDSA_SIGNATURE_376                                                               (32'h1118)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_377                                                           (32'h1003111c)
`define MLDSA_REG_MLDSA_SIGNATURE_377                                                               (32'h111c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_378                                                           (32'h10031120)
`define MLDSA_REG_MLDSA_SIGNATURE_378                                                               (32'h1120)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_379                                                           (32'h10031124)
`define MLDSA_REG_MLDSA_SIGNATURE_379                                                               (32'h1124)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_380                                                           (32'h10031128)
`define MLDSA_REG_MLDSA_SIGNATURE_380                                                               (32'h1128)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_381                                                           (32'h1003112c)
`define MLDSA_REG_MLDSA_SIGNATURE_381                                                               (32'h112c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_382                                                           (32'h10031130)
`define MLDSA_REG_MLDSA_SIGNATURE_382                                                               (32'h1130)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_383                                                           (32'h10031134)
`define MLDSA_REG_MLDSA_SIGNATURE_383                                                               (32'h1134)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_384                                                           (32'h10031138)
`define MLDSA_REG_MLDSA_SIGNATURE_384                                                               (32'h1138)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_385                                                           (32'h1003113c)
`define MLDSA_REG_MLDSA_SIGNATURE_385                                                               (32'h113c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_386                                                           (32'h10031140)
`define MLDSA_REG_MLDSA_SIGNATURE_386                                                               (32'h1140)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_387                                                           (32'h10031144)
`define MLDSA_REG_MLDSA_SIGNATURE_387                                                               (32'h1144)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_388                                                           (32'h10031148)
`define MLDSA_REG_MLDSA_SIGNATURE_388                                                               (32'h1148)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_389                                                           (32'h1003114c)
`define MLDSA_REG_MLDSA_SIGNATURE_389                                                               (32'h114c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_390                                                           (32'h10031150)
`define MLDSA_REG_MLDSA_SIGNATURE_390                                                               (32'h1150)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_391                                                           (32'h10031154)
`define MLDSA_REG_MLDSA_SIGNATURE_391                                                               (32'h1154)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_392                                                           (32'h10031158)
`define MLDSA_REG_MLDSA_SIGNATURE_392                                                               (32'h1158)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_393                                                           (32'h1003115c)
`define MLDSA_REG_MLDSA_SIGNATURE_393                                                               (32'h115c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_394                                                           (32'h10031160)
`define MLDSA_REG_MLDSA_SIGNATURE_394                                                               (32'h1160)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_395                                                           (32'h10031164)
`define MLDSA_REG_MLDSA_SIGNATURE_395                                                               (32'h1164)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_396                                                           (32'h10031168)
`define MLDSA_REG_MLDSA_SIGNATURE_396                                                               (32'h1168)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_397                                                           (32'h1003116c)
`define MLDSA_REG_MLDSA_SIGNATURE_397                                                               (32'h116c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_398                                                           (32'h10031170)
`define MLDSA_REG_MLDSA_SIGNATURE_398                                                               (32'h1170)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_399                                                           (32'h10031174)
`define MLDSA_REG_MLDSA_SIGNATURE_399                                                               (32'h1174)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_400                                                           (32'h10031178)
`define MLDSA_REG_MLDSA_SIGNATURE_400                                                               (32'h1178)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_401                                                           (32'h1003117c)
`define MLDSA_REG_MLDSA_SIGNATURE_401                                                               (32'h117c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_402                                                           (32'h10031180)
`define MLDSA_REG_MLDSA_SIGNATURE_402                                                               (32'h1180)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_403                                                           (32'h10031184)
`define MLDSA_REG_MLDSA_SIGNATURE_403                                                               (32'h1184)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_404                                                           (32'h10031188)
`define MLDSA_REG_MLDSA_SIGNATURE_404                                                               (32'h1188)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_405                                                           (32'h1003118c)
`define MLDSA_REG_MLDSA_SIGNATURE_405                                                               (32'h118c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_406                                                           (32'h10031190)
`define MLDSA_REG_MLDSA_SIGNATURE_406                                                               (32'h1190)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_407                                                           (32'h10031194)
`define MLDSA_REG_MLDSA_SIGNATURE_407                                                               (32'h1194)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_408                                                           (32'h10031198)
`define MLDSA_REG_MLDSA_SIGNATURE_408                                                               (32'h1198)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_409                                                           (32'h1003119c)
`define MLDSA_REG_MLDSA_SIGNATURE_409                                                               (32'h119c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_410                                                           (32'h100311a0)
`define MLDSA_REG_MLDSA_SIGNATURE_410                                                               (32'h11a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_411                                                           (32'h100311a4)
`define MLDSA_REG_MLDSA_SIGNATURE_411                                                               (32'h11a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_412                                                           (32'h100311a8)
`define MLDSA_REG_MLDSA_SIGNATURE_412                                                               (32'h11a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_413                                                           (32'h100311ac)
`define MLDSA_REG_MLDSA_SIGNATURE_413                                                               (32'h11ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_414                                                           (32'h100311b0)
`define MLDSA_REG_MLDSA_SIGNATURE_414                                                               (32'h11b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_415                                                           (32'h100311b4)
`define MLDSA_REG_MLDSA_SIGNATURE_415                                                               (32'h11b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_416                                                           (32'h100311b8)
`define MLDSA_REG_MLDSA_SIGNATURE_416                                                               (32'h11b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_417                                                           (32'h100311bc)
`define MLDSA_REG_MLDSA_SIGNATURE_417                                                               (32'h11bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_418                                                           (32'h100311c0)
`define MLDSA_REG_MLDSA_SIGNATURE_418                                                               (32'h11c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_419                                                           (32'h100311c4)
`define MLDSA_REG_MLDSA_SIGNATURE_419                                                               (32'h11c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_420                                                           (32'h100311c8)
`define MLDSA_REG_MLDSA_SIGNATURE_420                                                               (32'h11c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_421                                                           (32'h100311cc)
`define MLDSA_REG_MLDSA_SIGNATURE_421                                                               (32'h11cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_422                                                           (32'h100311d0)
`define MLDSA_REG_MLDSA_SIGNATURE_422                                                               (32'h11d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_423                                                           (32'h100311d4)
`define MLDSA_REG_MLDSA_SIGNATURE_423                                                               (32'h11d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_424                                                           (32'h100311d8)
`define MLDSA_REG_MLDSA_SIGNATURE_424                                                               (32'h11d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_425                                                           (32'h100311dc)
`define MLDSA_REG_MLDSA_SIGNATURE_425                                                               (32'h11dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_426                                                           (32'h100311e0)
`define MLDSA_REG_MLDSA_SIGNATURE_426                                                               (32'h11e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_427                                                           (32'h100311e4)
`define MLDSA_REG_MLDSA_SIGNATURE_427                                                               (32'h11e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_428                                                           (32'h100311e8)
`define MLDSA_REG_MLDSA_SIGNATURE_428                                                               (32'h11e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_429                                                           (32'h100311ec)
`define MLDSA_REG_MLDSA_SIGNATURE_429                                                               (32'h11ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_430                                                           (32'h100311f0)
`define MLDSA_REG_MLDSA_SIGNATURE_430                                                               (32'h11f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_431                                                           (32'h100311f4)
`define MLDSA_REG_MLDSA_SIGNATURE_431                                                               (32'h11f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_432                                                           (32'h100311f8)
`define MLDSA_REG_MLDSA_SIGNATURE_432                                                               (32'h11f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_433                                                           (32'h100311fc)
`define MLDSA_REG_MLDSA_SIGNATURE_433                                                               (32'h11fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_434                                                           (32'h10031200)
`define MLDSA_REG_MLDSA_SIGNATURE_434                                                               (32'h1200)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_435                                                           (32'h10031204)
`define MLDSA_REG_MLDSA_SIGNATURE_435                                                               (32'h1204)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_436                                                           (32'h10031208)
`define MLDSA_REG_MLDSA_SIGNATURE_436                                                               (32'h1208)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_437                                                           (32'h1003120c)
`define MLDSA_REG_MLDSA_SIGNATURE_437                                                               (32'h120c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_438                                                           (32'h10031210)
`define MLDSA_REG_MLDSA_SIGNATURE_438                                                               (32'h1210)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_439                                                           (32'h10031214)
`define MLDSA_REG_MLDSA_SIGNATURE_439                                                               (32'h1214)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_440                                                           (32'h10031218)
`define MLDSA_REG_MLDSA_SIGNATURE_440                                                               (32'h1218)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_441                                                           (32'h1003121c)
`define MLDSA_REG_MLDSA_SIGNATURE_441                                                               (32'h121c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_442                                                           (32'h10031220)
`define MLDSA_REG_MLDSA_SIGNATURE_442                                                               (32'h1220)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_443                                                           (32'h10031224)
`define MLDSA_REG_MLDSA_SIGNATURE_443                                                               (32'h1224)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_444                                                           (32'h10031228)
`define MLDSA_REG_MLDSA_SIGNATURE_444                                                               (32'h1228)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_445                                                           (32'h1003122c)
`define MLDSA_REG_MLDSA_SIGNATURE_445                                                               (32'h122c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_446                                                           (32'h10031230)
`define MLDSA_REG_MLDSA_SIGNATURE_446                                                               (32'h1230)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_447                                                           (32'h10031234)
`define MLDSA_REG_MLDSA_SIGNATURE_447                                                               (32'h1234)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_448                                                           (32'h10031238)
`define MLDSA_REG_MLDSA_SIGNATURE_448                                                               (32'h1238)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_449                                                           (32'h1003123c)
`define MLDSA_REG_MLDSA_SIGNATURE_449                                                               (32'h123c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_450                                                           (32'h10031240)
`define MLDSA_REG_MLDSA_SIGNATURE_450                                                               (32'h1240)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_451                                                           (32'h10031244)
`define MLDSA_REG_MLDSA_SIGNATURE_451                                                               (32'h1244)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_452                                                           (32'h10031248)
`define MLDSA_REG_MLDSA_SIGNATURE_452                                                               (32'h1248)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_453                                                           (32'h1003124c)
`define MLDSA_REG_MLDSA_SIGNATURE_453                                                               (32'h124c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_454                                                           (32'h10031250)
`define MLDSA_REG_MLDSA_SIGNATURE_454                                                               (32'h1250)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_455                                                           (32'h10031254)
`define MLDSA_REG_MLDSA_SIGNATURE_455                                                               (32'h1254)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_456                                                           (32'h10031258)
`define MLDSA_REG_MLDSA_SIGNATURE_456                                                               (32'h1258)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_457                                                           (32'h1003125c)
`define MLDSA_REG_MLDSA_SIGNATURE_457                                                               (32'h125c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_458                                                           (32'h10031260)
`define MLDSA_REG_MLDSA_SIGNATURE_458                                                               (32'h1260)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_459                                                           (32'h10031264)
`define MLDSA_REG_MLDSA_SIGNATURE_459                                                               (32'h1264)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_460                                                           (32'h10031268)
`define MLDSA_REG_MLDSA_SIGNATURE_460                                                               (32'h1268)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_461                                                           (32'h1003126c)
`define MLDSA_REG_MLDSA_SIGNATURE_461                                                               (32'h126c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_462                                                           (32'h10031270)
`define MLDSA_REG_MLDSA_SIGNATURE_462                                                               (32'h1270)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_463                                                           (32'h10031274)
`define MLDSA_REG_MLDSA_SIGNATURE_463                                                               (32'h1274)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_464                                                           (32'h10031278)
`define MLDSA_REG_MLDSA_SIGNATURE_464                                                               (32'h1278)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_465                                                           (32'h1003127c)
`define MLDSA_REG_MLDSA_SIGNATURE_465                                                               (32'h127c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_466                                                           (32'h10031280)
`define MLDSA_REG_MLDSA_SIGNATURE_466                                                               (32'h1280)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_467                                                           (32'h10031284)
`define MLDSA_REG_MLDSA_SIGNATURE_467                                                               (32'h1284)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_468                                                           (32'h10031288)
`define MLDSA_REG_MLDSA_SIGNATURE_468                                                               (32'h1288)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_469                                                           (32'h1003128c)
`define MLDSA_REG_MLDSA_SIGNATURE_469                                                               (32'h128c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_470                                                           (32'h10031290)
`define MLDSA_REG_MLDSA_SIGNATURE_470                                                               (32'h1290)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_471                                                           (32'h10031294)
`define MLDSA_REG_MLDSA_SIGNATURE_471                                                               (32'h1294)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_472                                                           (32'h10031298)
`define MLDSA_REG_MLDSA_SIGNATURE_472                                                               (32'h1298)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_473                                                           (32'h1003129c)
`define MLDSA_REG_MLDSA_SIGNATURE_473                                                               (32'h129c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_474                                                           (32'h100312a0)
`define MLDSA_REG_MLDSA_SIGNATURE_474                                                               (32'h12a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_475                                                           (32'h100312a4)
`define MLDSA_REG_MLDSA_SIGNATURE_475                                                               (32'h12a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_476                                                           (32'h100312a8)
`define MLDSA_REG_MLDSA_SIGNATURE_476                                                               (32'h12a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_477                                                           (32'h100312ac)
`define MLDSA_REG_MLDSA_SIGNATURE_477                                                               (32'h12ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_478                                                           (32'h100312b0)
`define MLDSA_REG_MLDSA_SIGNATURE_478                                                               (32'h12b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_479                                                           (32'h100312b4)
`define MLDSA_REG_MLDSA_SIGNATURE_479                                                               (32'h12b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_480                                                           (32'h100312b8)
`define MLDSA_REG_MLDSA_SIGNATURE_480                                                               (32'h12b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_481                                                           (32'h100312bc)
`define MLDSA_REG_MLDSA_SIGNATURE_481                                                               (32'h12bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_482                                                           (32'h100312c0)
`define MLDSA_REG_MLDSA_SIGNATURE_482                                                               (32'h12c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_483                                                           (32'h100312c4)
`define MLDSA_REG_MLDSA_SIGNATURE_483                                                               (32'h12c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_484                                                           (32'h100312c8)
`define MLDSA_REG_MLDSA_SIGNATURE_484                                                               (32'h12c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_485                                                           (32'h100312cc)
`define MLDSA_REG_MLDSA_SIGNATURE_485                                                               (32'h12cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_486                                                           (32'h100312d0)
`define MLDSA_REG_MLDSA_SIGNATURE_486                                                               (32'h12d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_487                                                           (32'h100312d4)
`define MLDSA_REG_MLDSA_SIGNATURE_487                                                               (32'h12d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_488                                                           (32'h100312d8)
`define MLDSA_REG_MLDSA_SIGNATURE_488                                                               (32'h12d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_489                                                           (32'h100312dc)
`define MLDSA_REG_MLDSA_SIGNATURE_489                                                               (32'h12dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_490                                                           (32'h100312e0)
`define MLDSA_REG_MLDSA_SIGNATURE_490                                                               (32'h12e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_491                                                           (32'h100312e4)
`define MLDSA_REG_MLDSA_SIGNATURE_491                                                               (32'h12e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_492                                                           (32'h100312e8)
`define MLDSA_REG_MLDSA_SIGNATURE_492                                                               (32'h12e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_493                                                           (32'h100312ec)
`define MLDSA_REG_MLDSA_SIGNATURE_493                                                               (32'h12ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_494                                                           (32'h100312f0)
`define MLDSA_REG_MLDSA_SIGNATURE_494                                                               (32'h12f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_495                                                           (32'h100312f4)
`define MLDSA_REG_MLDSA_SIGNATURE_495                                                               (32'h12f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_496                                                           (32'h100312f8)
`define MLDSA_REG_MLDSA_SIGNATURE_496                                                               (32'h12f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_497                                                           (32'h100312fc)
`define MLDSA_REG_MLDSA_SIGNATURE_497                                                               (32'h12fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_498                                                           (32'h10031300)
`define MLDSA_REG_MLDSA_SIGNATURE_498                                                               (32'h1300)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_499                                                           (32'h10031304)
`define MLDSA_REG_MLDSA_SIGNATURE_499                                                               (32'h1304)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_500                                                           (32'h10031308)
`define MLDSA_REG_MLDSA_SIGNATURE_500                                                               (32'h1308)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_501                                                           (32'h1003130c)
`define MLDSA_REG_MLDSA_SIGNATURE_501                                                               (32'h130c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_502                                                           (32'h10031310)
`define MLDSA_REG_MLDSA_SIGNATURE_502                                                               (32'h1310)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_503                                                           (32'h10031314)
`define MLDSA_REG_MLDSA_SIGNATURE_503                                                               (32'h1314)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_504                                                           (32'h10031318)
`define MLDSA_REG_MLDSA_SIGNATURE_504                                                               (32'h1318)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_505                                                           (32'h1003131c)
`define MLDSA_REG_MLDSA_SIGNATURE_505                                                               (32'h131c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_506                                                           (32'h10031320)
`define MLDSA_REG_MLDSA_SIGNATURE_506                                                               (32'h1320)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_507                                                           (32'h10031324)
`define MLDSA_REG_MLDSA_SIGNATURE_507                                                               (32'h1324)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_508                                                           (32'h10031328)
`define MLDSA_REG_MLDSA_SIGNATURE_508                                                               (32'h1328)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_509                                                           (32'h1003132c)
`define MLDSA_REG_MLDSA_SIGNATURE_509                                                               (32'h132c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_510                                                           (32'h10031330)
`define MLDSA_REG_MLDSA_SIGNATURE_510                                                               (32'h1330)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_511                                                           (32'h10031334)
`define MLDSA_REG_MLDSA_SIGNATURE_511                                                               (32'h1334)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_512                                                           (32'h10031338)
`define MLDSA_REG_MLDSA_SIGNATURE_512                                                               (32'h1338)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_513                                                           (32'h1003133c)
`define MLDSA_REG_MLDSA_SIGNATURE_513                                                               (32'h133c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_514                                                           (32'h10031340)
`define MLDSA_REG_MLDSA_SIGNATURE_514                                                               (32'h1340)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_515                                                           (32'h10031344)
`define MLDSA_REG_MLDSA_SIGNATURE_515                                                               (32'h1344)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_516                                                           (32'h10031348)
`define MLDSA_REG_MLDSA_SIGNATURE_516                                                               (32'h1348)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_517                                                           (32'h1003134c)
`define MLDSA_REG_MLDSA_SIGNATURE_517                                                               (32'h134c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_518                                                           (32'h10031350)
`define MLDSA_REG_MLDSA_SIGNATURE_518                                                               (32'h1350)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_519                                                           (32'h10031354)
`define MLDSA_REG_MLDSA_SIGNATURE_519                                                               (32'h1354)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_520                                                           (32'h10031358)
`define MLDSA_REG_MLDSA_SIGNATURE_520                                                               (32'h1358)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_521                                                           (32'h1003135c)
`define MLDSA_REG_MLDSA_SIGNATURE_521                                                               (32'h135c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_522                                                           (32'h10031360)
`define MLDSA_REG_MLDSA_SIGNATURE_522                                                               (32'h1360)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_523                                                           (32'h10031364)
`define MLDSA_REG_MLDSA_SIGNATURE_523                                                               (32'h1364)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_524                                                           (32'h10031368)
`define MLDSA_REG_MLDSA_SIGNATURE_524                                                               (32'h1368)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_525                                                           (32'h1003136c)
`define MLDSA_REG_MLDSA_SIGNATURE_525                                                               (32'h136c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_526                                                           (32'h10031370)
`define MLDSA_REG_MLDSA_SIGNATURE_526                                                               (32'h1370)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_527                                                           (32'h10031374)
`define MLDSA_REG_MLDSA_SIGNATURE_527                                                               (32'h1374)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_528                                                           (32'h10031378)
`define MLDSA_REG_MLDSA_SIGNATURE_528                                                               (32'h1378)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_529                                                           (32'h1003137c)
`define MLDSA_REG_MLDSA_SIGNATURE_529                                                               (32'h137c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_530                                                           (32'h10031380)
`define MLDSA_REG_MLDSA_SIGNATURE_530                                                               (32'h1380)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_531                                                           (32'h10031384)
`define MLDSA_REG_MLDSA_SIGNATURE_531                                                               (32'h1384)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_532                                                           (32'h10031388)
`define MLDSA_REG_MLDSA_SIGNATURE_532                                                               (32'h1388)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_533                                                           (32'h1003138c)
`define MLDSA_REG_MLDSA_SIGNATURE_533                                                               (32'h138c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_534                                                           (32'h10031390)
`define MLDSA_REG_MLDSA_SIGNATURE_534                                                               (32'h1390)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_535                                                           (32'h10031394)
`define MLDSA_REG_MLDSA_SIGNATURE_535                                                               (32'h1394)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_536                                                           (32'h10031398)
`define MLDSA_REG_MLDSA_SIGNATURE_536                                                               (32'h1398)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_537                                                           (32'h1003139c)
`define MLDSA_REG_MLDSA_SIGNATURE_537                                                               (32'h139c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_538                                                           (32'h100313a0)
`define MLDSA_REG_MLDSA_SIGNATURE_538                                                               (32'h13a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_539                                                           (32'h100313a4)
`define MLDSA_REG_MLDSA_SIGNATURE_539                                                               (32'h13a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_540                                                           (32'h100313a8)
`define MLDSA_REG_MLDSA_SIGNATURE_540                                                               (32'h13a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_541                                                           (32'h100313ac)
`define MLDSA_REG_MLDSA_SIGNATURE_541                                                               (32'h13ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_542                                                           (32'h100313b0)
`define MLDSA_REG_MLDSA_SIGNATURE_542                                                               (32'h13b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_543                                                           (32'h100313b4)
`define MLDSA_REG_MLDSA_SIGNATURE_543                                                               (32'h13b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_544                                                           (32'h100313b8)
`define MLDSA_REG_MLDSA_SIGNATURE_544                                                               (32'h13b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_545                                                           (32'h100313bc)
`define MLDSA_REG_MLDSA_SIGNATURE_545                                                               (32'h13bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_546                                                           (32'h100313c0)
`define MLDSA_REG_MLDSA_SIGNATURE_546                                                               (32'h13c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_547                                                           (32'h100313c4)
`define MLDSA_REG_MLDSA_SIGNATURE_547                                                               (32'h13c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_548                                                           (32'h100313c8)
`define MLDSA_REG_MLDSA_SIGNATURE_548                                                               (32'h13c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_549                                                           (32'h100313cc)
`define MLDSA_REG_MLDSA_SIGNATURE_549                                                               (32'h13cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_550                                                           (32'h100313d0)
`define MLDSA_REG_MLDSA_SIGNATURE_550                                                               (32'h13d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_551                                                           (32'h100313d4)
`define MLDSA_REG_MLDSA_SIGNATURE_551                                                               (32'h13d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_552                                                           (32'h100313d8)
`define MLDSA_REG_MLDSA_SIGNATURE_552                                                               (32'h13d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_553                                                           (32'h100313dc)
`define MLDSA_REG_MLDSA_SIGNATURE_553                                                               (32'h13dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_554                                                           (32'h100313e0)
`define MLDSA_REG_MLDSA_SIGNATURE_554                                                               (32'h13e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_555                                                           (32'h100313e4)
`define MLDSA_REG_MLDSA_SIGNATURE_555                                                               (32'h13e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_556                                                           (32'h100313e8)
`define MLDSA_REG_MLDSA_SIGNATURE_556                                                               (32'h13e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_557                                                           (32'h100313ec)
`define MLDSA_REG_MLDSA_SIGNATURE_557                                                               (32'h13ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_558                                                           (32'h100313f0)
`define MLDSA_REG_MLDSA_SIGNATURE_558                                                               (32'h13f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_559                                                           (32'h100313f4)
`define MLDSA_REG_MLDSA_SIGNATURE_559                                                               (32'h13f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_560                                                           (32'h100313f8)
`define MLDSA_REG_MLDSA_SIGNATURE_560                                                               (32'h13f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_561                                                           (32'h100313fc)
`define MLDSA_REG_MLDSA_SIGNATURE_561                                                               (32'h13fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_562                                                           (32'h10031400)
`define MLDSA_REG_MLDSA_SIGNATURE_562                                                               (32'h1400)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_563                                                           (32'h10031404)
`define MLDSA_REG_MLDSA_SIGNATURE_563                                                               (32'h1404)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_564                                                           (32'h10031408)
`define MLDSA_REG_MLDSA_SIGNATURE_564                                                               (32'h1408)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_565                                                           (32'h1003140c)
`define MLDSA_REG_MLDSA_SIGNATURE_565                                                               (32'h140c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_566                                                           (32'h10031410)
`define MLDSA_REG_MLDSA_SIGNATURE_566                                                               (32'h1410)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_567                                                           (32'h10031414)
`define MLDSA_REG_MLDSA_SIGNATURE_567                                                               (32'h1414)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_568                                                           (32'h10031418)
`define MLDSA_REG_MLDSA_SIGNATURE_568                                                               (32'h1418)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_569                                                           (32'h1003141c)
`define MLDSA_REG_MLDSA_SIGNATURE_569                                                               (32'h141c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_570                                                           (32'h10031420)
`define MLDSA_REG_MLDSA_SIGNATURE_570                                                               (32'h1420)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_571                                                           (32'h10031424)
`define MLDSA_REG_MLDSA_SIGNATURE_571                                                               (32'h1424)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_572                                                           (32'h10031428)
`define MLDSA_REG_MLDSA_SIGNATURE_572                                                               (32'h1428)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_573                                                           (32'h1003142c)
`define MLDSA_REG_MLDSA_SIGNATURE_573                                                               (32'h142c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_574                                                           (32'h10031430)
`define MLDSA_REG_MLDSA_SIGNATURE_574                                                               (32'h1430)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_575                                                           (32'h10031434)
`define MLDSA_REG_MLDSA_SIGNATURE_575                                                               (32'h1434)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_576                                                           (32'h10031438)
`define MLDSA_REG_MLDSA_SIGNATURE_576                                                               (32'h1438)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_577                                                           (32'h1003143c)
`define MLDSA_REG_MLDSA_SIGNATURE_577                                                               (32'h143c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_578                                                           (32'h10031440)
`define MLDSA_REG_MLDSA_SIGNATURE_578                                                               (32'h1440)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_579                                                           (32'h10031444)
`define MLDSA_REG_MLDSA_SIGNATURE_579                                                               (32'h1444)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_580                                                           (32'h10031448)
`define MLDSA_REG_MLDSA_SIGNATURE_580                                                               (32'h1448)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_581                                                           (32'h1003144c)
`define MLDSA_REG_MLDSA_SIGNATURE_581                                                               (32'h144c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_582                                                           (32'h10031450)
`define MLDSA_REG_MLDSA_SIGNATURE_582                                                               (32'h1450)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_583                                                           (32'h10031454)
`define MLDSA_REG_MLDSA_SIGNATURE_583                                                               (32'h1454)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_584                                                           (32'h10031458)
`define MLDSA_REG_MLDSA_SIGNATURE_584                                                               (32'h1458)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_585                                                           (32'h1003145c)
`define MLDSA_REG_MLDSA_SIGNATURE_585                                                               (32'h145c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_586                                                           (32'h10031460)
`define MLDSA_REG_MLDSA_SIGNATURE_586                                                               (32'h1460)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_587                                                           (32'h10031464)
`define MLDSA_REG_MLDSA_SIGNATURE_587                                                               (32'h1464)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_588                                                           (32'h10031468)
`define MLDSA_REG_MLDSA_SIGNATURE_588                                                               (32'h1468)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_589                                                           (32'h1003146c)
`define MLDSA_REG_MLDSA_SIGNATURE_589                                                               (32'h146c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_590                                                           (32'h10031470)
`define MLDSA_REG_MLDSA_SIGNATURE_590                                                               (32'h1470)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_591                                                           (32'h10031474)
`define MLDSA_REG_MLDSA_SIGNATURE_591                                                               (32'h1474)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_592                                                           (32'h10031478)
`define MLDSA_REG_MLDSA_SIGNATURE_592                                                               (32'h1478)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_593                                                           (32'h1003147c)
`define MLDSA_REG_MLDSA_SIGNATURE_593                                                               (32'h147c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_594                                                           (32'h10031480)
`define MLDSA_REG_MLDSA_SIGNATURE_594                                                               (32'h1480)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_595                                                           (32'h10031484)
`define MLDSA_REG_MLDSA_SIGNATURE_595                                                               (32'h1484)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_596                                                           (32'h10031488)
`define MLDSA_REG_MLDSA_SIGNATURE_596                                                               (32'h1488)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_597                                                           (32'h1003148c)
`define MLDSA_REG_MLDSA_SIGNATURE_597                                                               (32'h148c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_598                                                           (32'h10031490)
`define MLDSA_REG_MLDSA_SIGNATURE_598                                                               (32'h1490)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_599                                                           (32'h10031494)
`define MLDSA_REG_MLDSA_SIGNATURE_599                                                               (32'h1494)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_600                                                           (32'h10031498)
`define MLDSA_REG_MLDSA_SIGNATURE_600                                                               (32'h1498)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_601                                                           (32'h1003149c)
`define MLDSA_REG_MLDSA_SIGNATURE_601                                                               (32'h149c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_602                                                           (32'h100314a0)
`define MLDSA_REG_MLDSA_SIGNATURE_602                                                               (32'h14a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_603                                                           (32'h100314a4)
`define MLDSA_REG_MLDSA_SIGNATURE_603                                                               (32'h14a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_604                                                           (32'h100314a8)
`define MLDSA_REG_MLDSA_SIGNATURE_604                                                               (32'h14a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_605                                                           (32'h100314ac)
`define MLDSA_REG_MLDSA_SIGNATURE_605                                                               (32'h14ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_606                                                           (32'h100314b0)
`define MLDSA_REG_MLDSA_SIGNATURE_606                                                               (32'h14b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_607                                                           (32'h100314b4)
`define MLDSA_REG_MLDSA_SIGNATURE_607                                                               (32'h14b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_608                                                           (32'h100314b8)
`define MLDSA_REG_MLDSA_SIGNATURE_608                                                               (32'h14b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_609                                                           (32'h100314bc)
`define MLDSA_REG_MLDSA_SIGNATURE_609                                                               (32'h14bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_610                                                           (32'h100314c0)
`define MLDSA_REG_MLDSA_SIGNATURE_610                                                               (32'h14c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_611                                                           (32'h100314c4)
`define MLDSA_REG_MLDSA_SIGNATURE_611                                                               (32'h14c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_612                                                           (32'h100314c8)
`define MLDSA_REG_MLDSA_SIGNATURE_612                                                               (32'h14c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_613                                                           (32'h100314cc)
`define MLDSA_REG_MLDSA_SIGNATURE_613                                                               (32'h14cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_614                                                           (32'h100314d0)
`define MLDSA_REG_MLDSA_SIGNATURE_614                                                               (32'h14d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_615                                                           (32'h100314d4)
`define MLDSA_REG_MLDSA_SIGNATURE_615                                                               (32'h14d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_616                                                           (32'h100314d8)
`define MLDSA_REG_MLDSA_SIGNATURE_616                                                               (32'h14d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_617                                                           (32'h100314dc)
`define MLDSA_REG_MLDSA_SIGNATURE_617                                                               (32'h14dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_618                                                           (32'h100314e0)
`define MLDSA_REG_MLDSA_SIGNATURE_618                                                               (32'h14e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_619                                                           (32'h100314e4)
`define MLDSA_REG_MLDSA_SIGNATURE_619                                                               (32'h14e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_620                                                           (32'h100314e8)
`define MLDSA_REG_MLDSA_SIGNATURE_620                                                               (32'h14e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_621                                                           (32'h100314ec)
`define MLDSA_REG_MLDSA_SIGNATURE_621                                                               (32'h14ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_622                                                           (32'h100314f0)
`define MLDSA_REG_MLDSA_SIGNATURE_622                                                               (32'h14f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_623                                                           (32'h100314f4)
`define MLDSA_REG_MLDSA_SIGNATURE_623                                                               (32'h14f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_624                                                           (32'h100314f8)
`define MLDSA_REG_MLDSA_SIGNATURE_624                                                               (32'h14f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_625                                                           (32'h100314fc)
`define MLDSA_REG_MLDSA_SIGNATURE_625                                                               (32'h14fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_626                                                           (32'h10031500)
`define MLDSA_REG_MLDSA_SIGNATURE_626                                                               (32'h1500)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_627                                                           (32'h10031504)
`define MLDSA_REG_MLDSA_SIGNATURE_627                                                               (32'h1504)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_628                                                           (32'h10031508)
`define MLDSA_REG_MLDSA_SIGNATURE_628                                                               (32'h1508)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_629                                                           (32'h1003150c)
`define MLDSA_REG_MLDSA_SIGNATURE_629                                                               (32'h150c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_630                                                           (32'h10031510)
`define MLDSA_REG_MLDSA_SIGNATURE_630                                                               (32'h1510)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_631                                                           (32'h10031514)
`define MLDSA_REG_MLDSA_SIGNATURE_631                                                               (32'h1514)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_632                                                           (32'h10031518)
`define MLDSA_REG_MLDSA_SIGNATURE_632                                                               (32'h1518)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_633                                                           (32'h1003151c)
`define MLDSA_REG_MLDSA_SIGNATURE_633                                                               (32'h151c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_634                                                           (32'h10031520)
`define MLDSA_REG_MLDSA_SIGNATURE_634                                                               (32'h1520)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_635                                                           (32'h10031524)
`define MLDSA_REG_MLDSA_SIGNATURE_635                                                               (32'h1524)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_636                                                           (32'h10031528)
`define MLDSA_REG_MLDSA_SIGNATURE_636                                                               (32'h1528)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_637                                                           (32'h1003152c)
`define MLDSA_REG_MLDSA_SIGNATURE_637                                                               (32'h152c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_638                                                           (32'h10031530)
`define MLDSA_REG_MLDSA_SIGNATURE_638                                                               (32'h1530)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_639                                                           (32'h10031534)
`define MLDSA_REG_MLDSA_SIGNATURE_639                                                               (32'h1534)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_640                                                           (32'h10031538)
`define MLDSA_REG_MLDSA_SIGNATURE_640                                                               (32'h1538)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_641                                                           (32'h1003153c)
`define MLDSA_REG_MLDSA_SIGNATURE_641                                                               (32'h153c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_642                                                           (32'h10031540)
`define MLDSA_REG_MLDSA_SIGNATURE_642                                                               (32'h1540)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_643                                                           (32'h10031544)
`define MLDSA_REG_MLDSA_SIGNATURE_643                                                               (32'h1544)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_644                                                           (32'h10031548)
`define MLDSA_REG_MLDSA_SIGNATURE_644                                                               (32'h1548)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_645                                                           (32'h1003154c)
`define MLDSA_REG_MLDSA_SIGNATURE_645                                                               (32'h154c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_646                                                           (32'h10031550)
`define MLDSA_REG_MLDSA_SIGNATURE_646                                                               (32'h1550)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_647                                                           (32'h10031554)
`define MLDSA_REG_MLDSA_SIGNATURE_647                                                               (32'h1554)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_648                                                           (32'h10031558)
`define MLDSA_REG_MLDSA_SIGNATURE_648                                                               (32'h1558)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_649                                                           (32'h1003155c)
`define MLDSA_REG_MLDSA_SIGNATURE_649                                                               (32'h155c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_650                                                           (32'h10031560)
`define MLDSA_REG_MLDSA_SIGNATURE_650                                                               (32'h1560)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_651                                                           (32'h10031564)
`define MLDSA_REG_MLDSA_SIGNATURE_651                                                               (32'h1564)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_652                                                           (32'h10031568)
`define MLDSA_REG_MLDSA_SIGNATURE_652                                                               (32'h1568)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_653                                                           (32'h1003156c)
`define MLDSA_REG_MLDSA_SIGNATURE_653                                                               (32'h156c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_654                                                           (32'h10031570)
`define MLDSA_REG_MLDSA_SIGNATURE_654                                                               (32'h1570)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_655                                                           (32'h10031574)
`define MLDSA_REG_MLDSA_SIGNATURE_655                                                               (32'h1574)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_656                                                           (32'h10031578)
`define MLDSA_REG_MLDSA_SIGNATURE_656                                                               (32'h1578)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_657                                                           (32'h1003157c)
`define MLDSA_REG_MLDSA_SIGNATURE_657                                                               (32'h157c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_658                                                           (32'h10031580)
`define MLDSA_REG_MLDSA_SIGNATURE_658                                                               (32'h1580)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_659                                                           (32'h10031584)
`define MLDSA_REG_MLDSA_SIGNATURE_659                                                               (32'h1584)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_660                                                           (32'h10031588)
`define MLDSA_REG_MLDSA_SIGNATURE_660                                                               (32'h1588)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_661                                                           (32'h1003158c)
`define MLDSA_REG_MLDSA_SIGNATURE_661                                                               (32'h158c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_662                                                           (32'h10031590)
`define MLDSA_REG_MLDSA_SIGNATURE_662                                                               (32'h1590)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_663                                                           (32'h10031594)
`define MLDSA_REG_MLDSA_SIGNATURE_663                                                               (32'h1594)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_664                                                           (32'h10031598)
`define MLDSA_REG_MLDSA_SIGNATURE_664                                                               (32'h1598)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_665                                                           (32'h1003159c)
`define MLDSA_REG_MLDSA_SIGNATURE_665                                                               (32'h159c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_666                                                           (32'h100315a0)
`define MLDSA_REG_MLDSA_SIGNATURE_666                                                               (32'h15a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_667                                                           (32'h100315a4)
`define MLDSA_REG_MLDSA_SIGNATURE_667                                                               (32'h15a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_668                                                           (32'h100315a8)
`define MLDSA_REG_MLDSA_SIGNATURE_668                                                               (32'h15a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_669                                                           (32'h100315ac)
`define MLDSA_REG_MLDSA_SIGNATURE_669                                                               (32'h15ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_670                                                           (32'h100315b0)
`define MLDSA_REG_MLDSA_SIGNATURE_670                                                               (32'h15b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_671                                                           (32'h100315b4)
`define MLDSA_REG_MLDSA_SIGNATURE_671                                                               (32'h15b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_672                                                           (32'h100315b8)
`define MLDSA_REG_MLDSA_SIGNATURE_672                                                               (32'h15b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_673                                                           (32'h100315bc)
`define MLDSA_REG_MLDSA_SIGNATURE_673                                                               (32'h15bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_674                                                           (32'h100315c0)
`define MLDSA_REG_MLDSA_SIGNATURE_674                                                               (32'h15c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_675                                                           (32'h100315c4)
`define MLDSA_REG_MLDSA_SIGNATURE_675                                                               (32'h15c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_676                                                           (32'h100315c8)
`define MLDSA_REG_MLDSA_SIGNATURE_676                                                               (32'h15c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_677                                                           (32'h100315cc)
`define MLDSA_REG_MLDSA_SIGNATURE_677                                                               (32'h15cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_678                                                           (32'h100315d0)
`define MLDSA_REG_MLDSA_SIGNATURE_678                                                               (32'h15d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_679                                                           (32'h100315d4)
`define MLDSA_REG_MLDSA_SIGNATURE_679                                                               (32'h15d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_680                                                           (32'h100315d8)
`define MLDSA_REG_MLDSA_SIGNATURE_680                                                               (32'h15d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_681                                                           (32'h100315dc)
`define MLDSA_REG_MLDSA_SIGNATURE_681                                                               (32'h15dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_682                                                           (32'h100315e0)
`define MLDSA_REG_MLDSA_SIGNATURE_682                                                               (32'h15e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_683                                                           (32'h100315e4)
`define MLDSA_REG_MLDSA_SIGNATURE_683                                                               (32'h15e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_684                                                           (32'h100315e8)
`define MLDSA_REG_MLDSA_SIGNATURE_684                                                               (32'h15e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_685                                                           (32'h100315ec)
`define MLDSA_REG_MLDSA_SIGNATURE_685                                                               (32'h15ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_686                                                           (32'h100315f0)
`define MLDSA_REG_MLDSA_SIGNATURE_686                                                               (32'h15f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_687                                                           (32'h100315f4)
`define MLDSA_REG_MLDSA_SIGNATURE_687                                                               (32'h15f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_688                                                           (32'h100315f8)
`define MLDSA_REG_MLDSA_SIGNATURE_688                                                               (32'h15f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_689                                                           (32'h100315fc)
`define MLDSA_REG_MLDSA_SIGNATURE_689                                                               (32'h15fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_690                                                           (32'h10031600)
`define MLDSA_REG_MLDSA_SIGNATURE_690                                                               (32'h1600)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_691                                                           (32'h10031604)
`define MLDSA_REG_MLDSA_SIGNATURE_691                                                               (32'h1604)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_692                                                           (32'h10031608)
`define MLDSA_REG_MLDSA_SIGNATURE_692                                                               (32'h1608)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_693                                                           (32'h1003160c)
`define MLDSA_REG_MLDSA_SIGNATURE_693                                                               (32'h160c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_694                                                           (32'h10031610)
`define MLDSA_REG_MLDSA_SIGNATURE_694                                                               (32'h1610)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_695                                                           (32'h10031614)
`define MLDSA_REG_MLDSA_SIGNATURE_695                                                               (32'h1614)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_696                                                           (32'h10031618)
`define MLDSA_REG_MLDSA_SIGNATURE_696                                                               (32'h1618)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_697                                                           (32'h1003161c)
`define MLDSA_REG_MLDSA_SIGNATURE_697                                                               (32'h161c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_698                                                           (32'h10031620)
`define MLDSA_REG_MLDSA_SIGNATURE_698                                                               (32'h1620)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_699                                                           (32'h10031624)
`define MLDSA_REG_MLDSA_SIGNATURE_699                                                               (32'h1624)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_700                                                           (32'h10031628)
`define MLDSA_REG_MLDSA_SIGNATURE_700                                                               (32'h1628)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_701                                                           (32'h1003162c)
`define MLDSA_REG_MLDSA_SIGNATURE_701                                                               (32'h162c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_702                                                           (32'h10031630)
`define MLDSA_REG_MLDSA_SIGNATURE_702                                                               (32'h1630)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_703                                                           (32'h10031634)
`define MLDSA_REG_MLDSA_SIGNATURE_703                                                               (32'h1634)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_704                                                           (32'h10031638)
`define MLDSA_REG_MLDSA_SIGNATURE_704                                                               (32'h1638)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_705                                                           (32'h1003163c)
`define MLDSA_REG_MLDSA_SIGNATURE_705                                                               (32'h163c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_706                                                           (32'h10031640)
`define MLDSA_REG_MLDSA_SIGNATURE_706                                                               (32'h1640)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_707                                                           (32'h10031644)
`define MLDSA_REG_MLDSA_SIGNATURE_707                                                               (32'h1644)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_708                                                           (32'h10031648)
`define MLDSA_REG_MLDSA_SIGNATURE_708                                                               (32'h1648)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_709                                                           (32'h1003164c)
`define MLDSA_REG_MLDSA_SIGNATURE_709                                                               (32'h164c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_710                                                           (32'h10031650)
`define MLDSA_REG_MLDSA_SIGNATURE_710                                                               (32'h1650)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_711                                                           (32'h10031654)
`define MLDSA_REG_MLDSA_SIGNATURE_711                                                               (32'h1654)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_712                                                           (32'h10031658)
`define MLDSA_REG_MLDSA_SIGNATURE_712                                                               (32'h1658)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_713                                                           (32'h1003165c)
`define MLDSA_REG_MLDSA_SIGNATURE_713                                                               (32'h165c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_714                                                           (32'h10031660)
`define MLDSA_REG_MLDSA_SIGNATURE_714                                                               (32'h1660)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_715                                                           (32'h10031664)
`define MLDSA_REG_MLDSA_SIGNATURE_715                                                               (32'h1664)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_716                                                           (32'h10031668)
`define MLDSA_REG_MLDSA_SIGNATURE_716                                                               (32'h1668)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_717                                                           (32'h1003166c)
`define MLDSA_REG_MLDSA_SIGNATURE_717                                                               (32'h166c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_718                                                           (32'h10031670)
`define MLDSA_REG_MLDSA_SIGNATURE_718                                                               (32'h1670)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_719                                                           (32'h10031674)
`define MLDSA_REG_MLDSA_SIGNATURE_719                                                               (32'h1674)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_720                                                           (32'h10031678)
`define MLDSA_REG_MLDSA_SIGNATURE_720                                                               (32'h1678)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_721                                                           (32'h1003167c)
`define MLDSA_REG_MLDSA_SIGNATURE_721                                                               (32'h167c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_722                                                           (32'h10031680)
`define MLDSA_REG_MLDSA_SIGNATURE_722                                                               (32'h1680)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_723                                                           (32'h10031684)
`define MLDSA_REG_MLDSA_SIGNATURE_723                                                               (32'h1684)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_724                                                           (32'h10031688)
`define MLDSA_REG_MLDSA_SIGNATURE_724                                                               (32'h1688)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_725                                                           (32'h1003168c)
`define MLDSA_REG_MLDSA_SIGNATURE_725                                                               (32'h168c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_726                                                           (32'h10031690)
`define MLDSA_REG_MLDSA_SIGNATURE_726                                                               (32'h1690)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_727                                                           (32'h10031694)
`define MLDSA_REG_MLDSA_SIGNATURE_727                                                               (32'h1694)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_728                                                           (32'h10031698)
`define MLDSA_REG_MLDSA_SIGNATURE_728                                                               (32'h1698)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_729                                                           (32'h1003169c)
`define MLDSA_REG_MLDSA_SIGNATURE_729                                                               (32'h169c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_730                                                           (32'h100316a0)
`define MLDSA_REG_MLDSA_SIGNATURE_730                                                               (32'h16a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_731                                                           (32'h100316a4)
`define MLDSA_REG_MLDSA_SIGNATURE_731                                                               (32'h16a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_732                                                           (32'h100316a8)
`define MLDSA_REG_MLDSA_SIGNATURE_732                                                               (32'h16a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_733                                                           (32'h100316ac)
`define MLDSA_REG_MLDSA_SIGNATURE_733                                                               (32'h16ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_734                                                           (32'h100316b0)
`define MLDSA_REG_MLDSA_SIGNATURE_734                                                               (32'h16b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_735                                                           (32'h100316b4)
`define MLDSA_REG_MLDSA_SIGNATURE_735                                                               (32'h16b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_736                                                           (32'h100316b8)
`define MLDSA_REG_MLDSA_SIGNATURE_736                                                               (32'h16b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_737                                                           (32'h100316bc)
`define MLDSA_REG_MLDSA_SIGNATURE_737                                                               (32'h16bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_738                                                           (32'h100316c0)
`define MLDSA_REG_MLDSA_SIGNATURE_738                                                               (32'h16c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_739                                                           (32'h100316c4)
`define MLDSA_REG_MLDSA_SIGNATURE_739                                                               (32'h16c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_740                                                           (32'h100316c8)
`define MLDSA_REG_MLDSA_SIGNATURE_740                                                               (32'h16c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_741                                                           (32'h100316cc)
`define MLDSA_REG_MLDSA_SIGNATURE_741                                                               (32'h16cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_742                                                           (32'h100316d0)
`define MLDSA_REG_MLDSA_SIGNATURE_742                                                               (32'h16d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_743                                                           (32'h100316d4)
`define MLDSA_REG_MLDSA_SIGNATURE_743                                                               (32'h16d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_744                                                           (32'h100316d8)
`define MLDSA_REG_MLDSA_SIGNATURE_744                                                               (32'h16d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_745                                                           (32'h100316dc)
`define MLDSA_REG_MLDSA_SIGNATURE_745                                                               (32'h16dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_746                                                           (32'h100316e0)
`define MLDSA_REG_MLDSA_SIGNATURE_746                                                               (32'h16e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_747                                                           (32'h100316e4)
`define MLDSA_REG_MLDSA_SIGNATURE_747                                                               (32'h16e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_748                                                           (32'h100316e8)
`define MLDSA_REG_MLDSA_SIGNATURE_748                                                               (32'h16e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_749                                                           (32'h100316ec)
`define MLDSA_REG_MLDSA_SIGNATURE_749                                                               (32'h16ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_750                                                           (32'h100316f0)
`define MLDSA_REG_MLDSA_SIGNATURE_750                                                               (32'h16f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_751                                                           (32'h100316f4)
`define MLDSA_REG_MLDSA_SIGNATURE_751                                                               (32'h16f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_752                                                           (32'h100316f8)
`define MLDSA_REG_MLDSA_SIGNATURE_752                                                               (32'h16f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_753                                                           (32'h100316fc)
`define MLDSA_REG_MLDSA_SIGNATURE_753                                                               (32'h16fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_754                                                           (32'h10031700)
`define MLDSA_REG_MLDSA_SIGNATURE_754                                                               (32'h1700)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_755                                                           (32'h10031704)
`define MLDSA_REG_MLDSA_SIGNATURE_755                                                               (32'h1704)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_756                                                           (32'h10031708)
`define MLDSA_REG_MLDSA_SIGNATURE_756                                                               (32'h1708)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_757                                                           (32'h1003170c)
`define MLDSA_REG_MLDSA_SIGNATURE_757                                                               (32'h170c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_758                                                           (32'h10031710)
`define MLDSA_REG_MLDSA_SIGNATURE_758                                                               (32'h1710)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_759                                                           (32'h10031714)
`define MLDSA_REG_MLDSA_SIGNATURE_759                                                               (32'h1714)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_760                                                           (32'h10031718)
`define MLDSA_REG_MLDSA_SIGNATURE_760                                                               (32'h1718)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_761                                                           (32'h1003171c)
`define MLDSA_REG_MLDSA_SIGNATURE_761                                                               (32'h171c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_762                                                           (32'h10031720)
`define MLDSA_REG_MLDSA_SIGNATURE_762                                                               (32'h1720)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_763                                                           (32'h10031724)
`define MLDSA_REG_MLDSA_SIGNATURE_763                                                               (32'h1724)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_764                                                           (32'h10031728)
`define MLDSA_REG_MLDSA_SIGNATURE_764                                                               (32'h1728)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_765                                                           (32'h1003172c)
`define MLDSA_REG_MLDSA_SIGNATURE_765                                                               (32'h172c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_766                                                           (32'h10031730)
`define MLDSA_REG_MLDSA_SIGNATURE_766                                                               (32'h1730)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_767                                                           (32'h10031734)
`define MLDSA_REG_MLDSA_SIGNATURE_767                                                               (32'h1734)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_768                                                           (32'h10031738)
`define MLDSA_REG_MLDSA_SIGNATURE_768                                                               (32'h1738)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_769                                                           (32'h1003173c)
`define MLDSA_REG_MLDSA_SIGNATURE_769                                                               (32'h173c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_770                                                           (32'h10031740)
`define MLDSA_REG_MLDSA_SIGNATURE_770                                                               (32'h1740)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_771                                                           (32'h10031744)
`define MLDSA_REG_MLDSA_SIGNATURE_771                                                               (32'h1744)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_772                                                           (32'h10031748)
`define MLDSA_REG_MLDSA_SIGNATURE_772                                                               (32'h1748)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_773                                                           (32'h1003174c)
`define MLDSA_REG_MLDSA_SIGNATURE_773                                                               (32'h174c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_774                                                           (32'h10031750)
`define MLDSA_REG_MLDSA_SIGNATURE_774                                                               (32'h1750)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_775                                                           (32'h10031754)
`define MLDSA_REG_MLDSA_SIGNATURE_775                                                               (32'h1754)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_776                                                           (32'h10031758)
`define MLDSA_REG_MLDSA_SIGNATURE_776                                                               (32'h1758)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_777                                                           (32'h1003175c)
`define MLDSA_REG_MLDSA_SIGNATURE_777                                                               (32'h175c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_778                                                           (32'h10031760)
`define MLDSA_REG_MLDSA_SIGNATURE_778                                                               (32'h1760)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_779                                                           (32'h10031764)
`define MLDSA_REG_MLDSA_SIGNATURE_779                                                               (32'h1764)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_780                                                           (32'h10031768)
`define MLDSA_REG_MLDSA_SIGNATURE_780                                                               (32'h1768)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_781                                                           (32'h1003176c)
`define MLDSA_REG_MLDSA_SIGNATURE_781                                                               (32'h176c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_782                                                           (32'h10031770)
`define MLDSA_REG_MLDSA_SIGNATURE_782                                                               (32'h1770)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_783                                                           (32'h10031774)
`define MLDSA_REG_MLDSA_SIGNATURE_783                                                               (32'h1774)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_784                                                           (32'h10031778)
`define MLDSA_REG_MLDSA_SIGNATURE_784                                                               (32'h1778)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_785                                                           (32'h1003177c)
`define MLDSA_REG_MLDSA_SIGNATURE_785                                                               (32'h177c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_786                                                           (32'h10031780)
`define MLDSA_REG_MLDSA_SIGNATURE_786                                                               (32'h1780)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_787                                                           (32'h10031784)
`define MLDSA_REG_MLDSA_SIGNATURE_787                                                               (32'h1784)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_788                                                           (32'h10031788)
`define MLDSA_REG_MLDSA_SIGNATURE_788                                                               (32'h1788)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_789                                                           (32'h1003178c)
`define MLDSA_REG_MLDSA_SIGNATURE_789                                                               (32'h178c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_790                                                           (32'h10031790)
`define MLDSA_REG_MLDSA_SIGNATURE_790                                                               (32'h1790)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_791                                                           (32'h10031794)
`define MLDSA_REG_MLDSA_SIGNATURE_791                                                               (32'h1794)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_792                                                           (32'h10031798)
`define MLDSA_REG_MLDSA_SIGNATURE_792                                                               (32'h1798)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_793                                                           (32'h1003179c)
`define MLDSA_REG_MLDSA_SIGNATURE_793                                                               (32'h179c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_794                                                           (32'h100317a0)
`define MLDSA_REG_MLDSA_SIGNATURE_794                                                               (32'h17a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_795                                                           (32'h100317a4)
`define MLDSA_REG_MLDSA_SIGNATURE_795                                                               (32'h17a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_796                                                           (32'h100317a8)
`define MLDSA_REG_MLDSA_SIGNATURE_796                                                               (32'h17a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_797                                                           (32'h100317ac)
`define MLDSA_REG_MLDSA_SIGNATURE_797                                                               (32'h17ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_798                                                           (32'h100317b0)
`define MLDSA_REG_MLDSA_SIGNATURE_798                                                               (32'h17b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_799                                                           (32'h100317b4)
`define MLDSA_REG_MLDSA_SIGNATURE_799                                                               (32'h17b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_800                                                           (32'h100317b8)
`define MLDSA_REG_MLDSA_SIGNATURE_800                                                               (32'h17b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_801                                                           (32'h100317bc)
`define MLDSA_REG_MLDSA_SIGNATURE_801                                                               (32'h17bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_802                                                           (32'h100317c0)
`define MLDSA_REG_MLDSA_SIGNATURE_802                                                               (32'h17c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_803                                                           (32'h100317c4)
`define MLDSA_REG_MLDSA_SIGNATURE_803                                                               (32'h17c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_804                                                           (32'h100317c8)
`define MLDSA_REG_MLDSA_SIGNATURE_804                                                               (32'h17c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_805                                                           (32'h100317cc)
`define MLDSA_REG_MLDSA_SIGNATURE_805                                                               (32'h17cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_806                                                           (32'h100317d0)
`define MLDSA_REG_MLDSA_SIGNATURE_806                                                               (32'h17d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_807                                                           (32'h100317d4)
`define MLDSA_REG_MLDSA_SIGNATURE_807                                                               (32'h17d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_808                                                           (32'h100317d8)
`define MLDSA_REG_MLDSA_SIGNATURE_808                                                               (32'h17d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_809                                                           (32'h100317dc)
`define MLDSA_REG_MLDSA_SIGNATURE_809                                                               (32'h17dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_810                                                           (32'h100317e0)
`define MLDSA_REG_MLDSA_SIGNATURE_810                                                               (32'h17e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_811                                                           (32'h100317e4)
`define MLDSA_REG_MLDSA_SIGNATURE_811                                                               (32'h17e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_812                                                           (32'h100317e8)
`define MLDSA_REG_MLDSA_SIGNATURE_812                                                               (32'h17e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_813                                                           (32'h100317ec)
`define MLDSA_REG_MLDSA_SIGNATURE_813                                                               (32'h17ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_814                                                           (32'h100317f0)
`define MLDSA_REG_MLDSA_SIGNATURE_814                                                               (32'h17f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_815                                                           (32'h100317f4)
`define MLDSA_REG_MLDSA_SIGNATURE_815                                                               (32'h17f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_816                                                           (32'h100317f8)
`define MLDSA_REG_MLDSA_SIGNATURE_816                                                               (32'h17f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_817                                                           (32'h100317fc)
`define MLDSA_REG_MLDSA_SIGNATURE_817                                                               (32'h17fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_818                                                           (32'h10031800)
`define MLDSA_REG_MLDSA_SIGNATURE_818                                                               (32'h1800)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_819                                                           (32'h10031804)
`define MLDSA_REG_MLDSA_SIGNATURE_819                                                               (32'h1804)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_820                                                           (32'h10031808)
`define MLDSA_REG_MLDSA_SIGNATURE_820                                                               (32'h1808)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_821                                                           (32'h1003180c)
`define MLDSA_REG_MLDSA_SIGNATURE_821                                                               (32'h180c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_822                                                           (32'h10031810)
`define MLDSA_REG_MLDSA_SIGNATURE_822                                                               (32'h1810)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_823                                                           (32'h10031814)
`define MLDSA_REG_MLDSA_SIGNATURE_823                                                               (32'h1814)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_824                                                           (32'h10031818)
`define MLDSA_REG_MLDSA_SIGNATURE_824                                                               (32'h1818)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_825                                                           (32'h1003181c)
`define MLDSA_REG_MLDSA_SIGNATURE_825                                                               (32'h181c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_826                                                           (32'h10031820)
`define MLDSA_REG_MLDSA_SIGNATURE_826                                                               (32'h1820)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_827                                                           (32'h10031824)
`define MLDSA_REG_MLDSA_SIGNATURE_827                                                               (32'h1824)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_828                                                           (32'h10031828)
`define MLDSA_REG_MLDSA_SIGNATURE_828                                                               (32'h1828)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_829                                                           (32'h1003182c)
`define MLDSA_REG_MLDSA_SIGNATURE_829                                                               (32'h182c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_830                                                           (32'h10031830)
`define MLDSA_REG_MLDSA_SIGNATURE_830                                                               (32'h1830)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_831                                                           (32'h10031834)
`define MLDSA_REG_MLDSA_SIGNATURE_831                                                               (32'h1834)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_832                                                           (32'h10031838)
`define MLDSA_REG_MLDSA_SIGNATURE_832                                                               (32'h1838)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_833                                                           (32'h1003183c)
`define MLDSA_REG_MLDSA_SIGNATURE_833                                                               (32'h183c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_834                                                           (32'h10031840)
`define MLDSA_REG_MLDSA_SIGNATURE_834                                                               (32'h1840)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_835                                                           (32'h10031844)
`define MLDSA_REG_MLDSA_SIGNATURE_835                                                               (32'h1844)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_836                                                           (32'h10031848)
`define MLDSA_REG_MLDSA_SIGNATURE_836                                                               (32'h1848)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_837                                                           (32'h1003184c)
`define MLDSA_REG_MLDSA_SIGNATURE_837                                                               (32'h184c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_838                                                           (32'h10031850)
`define MLDSA_REG_MLDSA_SIGNATURE_838                                                               (32'h1850)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_839                                                           (32'h10031854)
`define MLDSA_REG_MLDSA_SIGNATURE_839                                                               (32'h1854)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_840                                                           (32'h10031858)
`define MLDSA_REG_MLDSA_SIGNATURE_840                                                               (32'h1858)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_841                                                           (32'h1003185c)
`define MLDSA_REG_MLDSA_SIGNATURE_841                                                               (32'h185c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_842                                                           (32'h10031860)
`define MLDSA_REG_MLDSA_SIGNATURE_842                                                               (32'h1860)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_843                                                           (32'h10031864)
`define MLDSA_REG_MLDSA_SIGNATURE_843                                                               (32'h1864)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_844                                                           (32'h10031868)
`define MLDSA_REG_MLDSA_SIGNATURE_844                                                               (32'h1868)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_845                                                           (32'h1003186c)
`define MLDSA_REG_MLDSA_SIGNATURE_845                                                               (32'h186c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_846                                                           (32'h10031870)
`define MLDSA_REG_MLDSA_SIGNATURE_846                                                               (32'h1870)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_847                                                           (32'h10031874)
`define MLDSA_REG_MLDSA_SIGNATURE_847                                                               (32'h1874)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_848                                                           (32'h10031878)
`define MLDSA_REG_MLDSA_SIGNATURE_848                                                               (32'h1878)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_849                                                           (32'h1003187c)
`define MLDSA_REG_MLDSA_SIGNATURE_849                                                               (32'h187c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_850                                                           (32'h10031880)
`define MLDSA_REG_MLDSA_SIGNATURE_850                                                               (32'h1880)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_851                                                           (32'h10031884)
`define MLDSA_REG_MLDSA_SIGNATURE_851                                                               (32'h1884)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_852                                                           (32'h10031888)
`define MLDSA_REG_MLDSA_SIGNATURE_852                                                               (32'h1888)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_853                                                           (32'h1003188c)
`define MLDSA_REG_MLDSA_SIGNATURE_853                                                               (32'h188c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_854                                                           (32'h10031890)
`define MLDSA_REG_MLDSA_SIGNATURE_854                                                               (32'h1890)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_855                                                           (32'h10031894)
`define MLDSA_REG_MLDSA_SIGNATURE_855                                                               (32'h1894)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_856                                                           (32'h10031898)
`define MLDSA_REG_MLDSA_SIGNATURE_856                                                               (32'h1898)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_857                                                           (32'h1003189c)
`define MLDSA_REG_MLDSA_SIGNATURE_857                                                               (32'h189c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_858                                                           (32'h100318a0)
`define MLDSA_REG_MLDSA_SIGNATURE_858                                                               (32'h18a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_859                                                           (32'h100318a4)
`define MLDSA_REG_MLDSA_SIGNATURE_859                                                               (32'h18a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_860                                                           (32'h100318a8)
`define MLDSA_REG_MLDSA_SIGNATURE_860                                                               (32'h18a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_861                                                           (32'h100318ac)
`define MLDSA_REG_MLDSA_SIGNATURE_861                                                               (32'h18ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_862                                                           (32'h100318b0)
`define MLDSA_REG_MLDSA_SIGNATURE_862                                                               (32'h18b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_863                                                           (32'h100318b4)
`define MLDSA_REG_MLDSA_SIGNATURE_863                                                               (32'h18b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_864                                                           (32'h100318b8)
`define MLDSA_REG_MLDSA_SIGNATURE_864                                                               (32'h18b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_865                                                           (32'h100318bc)
`define MLDSA_REG_MLDSA_SIGNATURE_865                                                               (32'h18bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_866                                                           (32'h100318c0)
`define MLDSA_REG_MLDSA_SIGNATURE_866                                                               (32'h18c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_867                                                           (32'h100318c4)
`define MLDSA_REG_MLDSA_SIGNATURE_867                                                               (32'h18c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_868                                                           (32'h100318c8)
`define MLDSA_REG_MLDSA_SIGNATURE_868                                                               (32'h18c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_869                                                           (32'h100318cc)
`define MLDSA_REG_MLDSA_SIGNATURE_869                                                               (32'h18cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_870                                                           (32'h100318d0)
`define MLDSA_REG_MLDSA_SIGNATURE_870                                                               (32'h18d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_871                                                           (32'h100318d4)
`define MLDSA_REG_MLDSA_SIGNATURE_871                                                               (32'h18d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_872                                                           (32'h100318d8)
`define MLDSA_REG_MLDSA_SIGNATURE_872                                                               (32'h18d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_873                                                           (32'h100318dc)
`define MLDSA_REG_MLDSA_SIGNATURE_873                                                               (32'h18dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_874                                                           (32'h100318e0)
`define MLDSA_REG_MLDSA_SIGNATURE_874                                                               (32'h18e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_875                                                           (32'h100318e4)
`define MLDSA_REG_MLDSA_SIGNATURE_875                                                               (32'h18e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_876                                                           (32'h100318e8)
`define MLDSA_REG_MLDSA_SIGNATURE_876                                                               (32'h18e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_877                                                           (32'h100318ec)
`define MLDSA_REG_MLDSA_SIGNATURE_877                                                               (32'h18ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_878                                                           (32'h100318f0)
`define MLDSA_REG_MLDSA_SIGNATURE_878                                                               (32'h18f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_879                                                           (32'h100318f4)
`define MLDSA_REG_MLDSA_SIGNATURE_879                                                               (32'h18f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_880                                                           (32'h100318f8)
`define MLDSA_REG_MLDSA_SIGNATURE_880                                                               (32'h18f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_881                                                           (32'h100318fc)
`define MLDSA_REG_MLDSA_SIGNATURE_881                                                               (32'h18fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_882                                                           (32'h10031900)
`define MLDSA_REG_MLDSA_SIGNATURE_882                                                               (32'h1900)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_883                                                           (32'h10031904)
`define MLDSA_REG_MLDSA_SIGNATURE_883                                                               (32'h1904)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_884                                                           (32'h10031908)
`define MLDSA_REG_MLDSA_SIGNATURE_884                                                               (32'h1908)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_885                                                           (32'h1003190c)
`define MLDSA_REG_MLDSA_SIGNATURE_885                                                               (32'h190c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_886                                                           (32'h10031910)
`define MLDSA_REG_MLDSA_SIGNATURE_886                                                               (32'h1910)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_887                                                           (32'h10031914)
`define MLDSA_REG_MLDSA_SIGNATURE_887                                                               (32'h1914)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_888                                                           (32'h10031918)
`define MLDSA_REG_MLDSA_SIGNATURE_888                                                               (32'h1918)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_889                                                           (32'h1003191c)
`define MLDSA_REG_MLDSA_SIGNATURE_889                                                               (32'h191c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_890                                                           (32'h10031920)
`define MLDSA_REG_MLDSA_SIGNATURE_890                                                               (32'h1920)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_891                                                           (32'h10031924)
`define MLDSA_REG_MLDSA_SIGNATURE_891                                                               (32'h1924)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_892                                                           (32'h10031928)
`define MLDSA_REG_MLDSA_SIGNATURE_892                                                               (32'h1928)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_893                                                           (32'h1003192c)
`define MLDSA_REG_MLDSA_SIGNATURE_893                                                               (32'h192c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_894                                                           (32'h10031930)
`define MLDSA_REG_MLDSA_SIGNATURE_894                                                               (32'h1930)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_895                                                           (32'h10031934)
`define MLDSA_REG_MLDSA_SIGNATURE_895                                                               (32'h1934)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_896                                                           (32'h10031938)
`define MLDSA_REG_MLDSA_SIGNATURE_896                                                               (32'h1938)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_897                                                           (32'h1003193c)
`define MLDSA_REG_MLDSA_SIGNATURE_897                                                               (32'h193c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_898                                                           (32'h10031940)
`define MLDSA_REG_MLDSA_SIGNATURE_898                                                               (32'h1940)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_899                                                           (32'h10031944)
`define MLDSA_REG_MLDSA_SIGNATURE_899                                                               (32'h1944)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_900                                                           (32'h10031948)
`define MLDSA_REG_MLDSA_SIGNATURE_900                                                               (32'h1948)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_901                                                           (32'h1003194c)
`define MLDSA_REG_MLDSA_SIGNATURE_901                                                               (32'h194c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_902                                                           (32'h10031950)
`define MLDSA_REG_MLDSA_SIGNATURE_902                                                               (32'h1950)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_903                                                           (32'h10031954)
`define MLDSA_REG_MLDSA_SIGNATURE_903                                                               (32'h1954)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_904                                                           (32'h10031958)
`define MLDSA_REG_MLDSA_SIGNATURE_904                                                               (32'h1958)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_905                                                           (32'h1003195c)
`define MLDSA_REG_MLDSA_SIGNATURE_905                                                               (32'h195c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_906                                                           (32'h10031960)
`define MLDSA_REG_MLDSA_SIGNATURE_906                                                               (32'h1960)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_907                                                           (32'h10031964)
`define MLDSA_REG_MLDSA_SIGNATURE_907                                                               (32'h1964)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_908                                                           (32'h10031968)
`define MLDSA_REG_MLDSA_SIGNATURE_908                                                               (32'h1968)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_909                                                           (32'h1003196c)
`define MLDSA_REG_MLDSA_SIGNATURE_909                                                               (32'h196c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_910                                                           (32'h10031970)
`define MLDSA_REG_MLDSA_SIGNATURE_910                                                               (32'h1970)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_911                                                           (32'h10031974)
`define MLDSA_REG_MLDSA_SIGNATURE_911                                                               (32'h1974)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_912                                                           (32'h10031978)
`define MLDSA_REG_MLDSA_SIGNATURE_912                                                               (32'h1978)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_913                                                           (32'h1003197c)
`define MLDSA_REG_MLDSA_SIGNATURE_913                                                               (32'h197c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_914                                                           (32'h10031980)
`define MLDSA_REG_MLDSA_SIGNATURE_914                                                               (32'h1980)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_915                                                           (32'h10031984)
`define MLDSA_REG_MLDSA_SIGNATURE_915                                                               (32'h1984)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_916                                                           (32'h10031988)
`define MLDSA_REG_MLDSA_SIGNATURE_916                                                               (32'h1988)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_917                                                           (32'h1003198c)
`define MLDSA_REG_MLDSA_SIGNATURE_917                                                               (32'h198c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_918                                                           (32'h10031990)
`define MLDSA_REG_MLDSA_SIGNATURE_918                                                               (32'h1990)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_919                                                           (32'h10031994)
`define MLDSA_REG_MLDSA_SIGNATURE_919                                                               (32'h1994)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_920                                                           (32'h10031998)
`define MLDSA_REG_MLDSA_SIGNATURE_920                                                               (32'h1998)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_921                                                           (32'h1003199c)
`define MLDSA_REG_MLDSA_SIGNATURE_921                                                               (32'h199c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_922                                                           (32'h100319a0)
`define MLDSA_REG_MLDSA_SIGNATURE_922                                                               (32'h19a0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_923                                                           (32'h100319a4)
`define MLDSA_REG_MLDSA_SIGNATURE_923                                                               (32'h19a4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_924                                                           (32'h100319a8)
`define MLDSA_REG_MLDSA_SIGNATURE_924                                                               (32'h19a8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_925                                                           (32'h100319ac)
`define MLDSA_REG_MLDSA_SIGNATURE_925                                                               (32'h19ac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_926                                                           (32'h100319b0)
`define MLDSA_REG_MLDSA_SIGNATURE_926                                                               (32'h19b0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_927                                                           (32'h100319b4)
`define MLDSA_REG_MLDSA_SIGNATURE_927                                                               (32'h19b4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_928                                                           (32'h100319b8)
`define MLDSA_REG_MLDSA_SIGNATURE_928                                                               (32'h19b8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_929                                                           (32'h100319bc)
`define MLDSA_REG_MLDSA_SIGNATURE_929                                                               (32'h19bc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_930                                                           (32'h100319c0)
`define MLDSA_REG_MLDSA_SIGNATURE_930                                                               (32'h19c0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_931                                                           (32'h100319c4)
`define MLDSA_REG_MLDSA_SIGNATURE_931                                                               (32'h19c4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_932                                                           (32'h100319c8)
`define MLDSA_REG_MLDSA_SIGNATURE_932                                                               (32'h19c8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_933                                                           (32'h100319cc)
`define MLDSA_REG_MLDSA_SIGNATURE_933                                                               (32'h19cc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_934                                                           (32'h100319d0)
`define MLDSA_REG_MLDSA_SIGNATURE_934                                                               (32'h19d0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_935                                                           (32'h100319d4)
`define MLDSA_REG_MLDSA_SIGNATURE_935                                                               (32'h19d4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_936                                                           (32'h100319d8)
`define MLDSA_REG_MLDSA_SIGNATURE_936                                                               (32'h19d8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_937                                                           (32'h100319dc)
`define MLDSA_REG_MLDSA_SIGNATURE_937                                                               (32'h19dc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_938                                                           (32'h100319e0)
`define MLDSA_REG_MLDSA_SIGNATURE_938                                                               (32'h19e0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_939                                                           (32'h100319e4)
`define MLDSA_REG_MLDSA_SIGNATURE_939                                                               (32'h19e4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_940                                                           (32'h100319e8)
`define MLDSA_REG_MLDSA_SIGNATURE_940                                                               (32'h19e8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_941                                                           (32'h100319ec)
`define MLDSA_REG_MLDSA_SIGNATURE_941                                                               (32'h19ec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_942                                                           (32'h100319f0)
`define MLDSA_REG_MLDSA_SIGNATURE_942                                                               (32'h19f0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_943                                                           (32'h100319f4)
`define MLDSA_REG_MLDSA_SIGNATURE_943                                                               (32'h19f4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_944                                                           (32'h100319f8)
`define MLDSA_REG_MLDSA_SIGNATURE_944                                                               (32'h19f8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_945                                                           (32'h100319fc)
`define MLDSA_REG_MLDSA_SIGNATURE_945                                                               (32'h19fc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_946                                                           (32'h10031a00)
`define MLDSA_REG_MLDSA_SIGNATURE_946                                                               (32'h1a00)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_947                                                           (32'h10031a04)
`define MLDSA_REG_MLDSA_SIGNATURE_947                                                               (32'h1a04)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_948                                                           (32'h10031a08)
`define MLDSA_REG_MLDSA_SIGNATURE_948                                                               (32'h1a08)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_949                                                           (32'h10031a0c)
`define MLDSA_REG_MLDSA_SIGNATURE_949                                                               (32'h1a0c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_950                                                           (32'h10031a10)
`define MLDSA_REG_MLDSA_SIGNATURE_950                                                               (32'h1a10)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_951                                                           (32'h10031a14)
`define MLDSA_REG_MLDSA_SIGNATURE_951                                                               (32'h1a14)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_952                                                           (32'h10031a18)
`define MLDSA_REG_MLDSA_SIGNATURE_952                                                               (32'h1a18)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_953                                                           (32'h10031a1c)
`define MLDSA_REG_MLDSA_SIGNATURE_953                                                               (32'h1a1c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_954                                                           (32'h10031a20)
`define MLDSA_REG_MLDSA_SIGNATURE_954                                                               (32'h1a20)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_955                                                           (32'h10031a24)
`define MLDSA_REG_MLDSA_SIGNATURE_955                                                               (32'h1a24)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_956                                                           (32'h10031a28)
`define MLDSA_REG_MLDSA_SIGNATURE_956                                                               (32'h1a28)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_957                                                           (32'h10031a2c)
`define MLDSA_REG_MLDSA_SIGNATURE_957                                                               (32'h1a2c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_958                                                           (32'h10031a30)
`define MLDSA_REG_MLDSA_SIGNATURE_958                                                               (32'h1a30)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_959                                                           (32'h10031a34)
`define MLDSA_REG_MLDSA_SIGNATURE_959                                                               (32'h1a34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_960                                                           (32'h10031a38)
`define MLDSA_REG_MLDSA_SIGNATURE_960                                                               (32'h1a38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_961                                                           (32'h10031a3c)
`define MLDSA_REG_MLDSA_SIGNATURE_961                                                               (32'h1a3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_962                                                           (32'h10031a40)
`define MLDSA_REG_MLDSA_SIGNATURE_962                                                               (32'h1a40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_963                                                           (32'h10031a44)
`define MLDSA_REG_MLDSA_SIGNATURE_963                                                               (32'h1a44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_964                                                           (32'h10031a48)
`define MLDSA_REG_MLDSA_SIGNATURE_964                                                               (32'h1a48)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_965                                                           (32'h10031a4c)
`define MLDSA_REG_MLDSA_SIGNATURE_965                                                               (32'h1a4c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_966                                                           (32'h10031a50)
`define MLDSA_REG_MLDSA_SIGNATURE_966                                                               (32'h1a50)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_967                                                           (32'h10031a54)
`define MLDSA_REG_MLDSA_SIGNATURE_967                                                               (32'h1a54)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_968                                                           (32'h10031a58)
`define MLDSA_REG_MLDSA_SIGNATURE_968                                                               (32'h1a58)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_969                                                           (32'h10031a5c)
`define MLDSA_REG_MLDSA_SIGNATURE_969                                                               (32'h1a5c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_970                                                           (32'h10031a60)
`define MLDSA_REG_MLDSA_SIGNATURE_970                                                               (32'h1a60)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_971                                                           (32'h10031a64)
`define MLDSA_REG_MLDSA_SIGNATURE_971                                                               (32'h1a64)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_972                                                           (32'h10031a68)
`define MLDSA_REG_MLDSA_SIGNATURE_972                                                               (32'h1a68)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_973                                                           (32'h10031a6c)
`define MLDSA_REG_MLDSA_SIGNATURE_973                                                               (32'h1a6c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_974                                                           (32'h10031a70)
`define MLDSA_REG_MLDSA_SIGNATURE_974                                                               (32'h1a70)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_975                                                           (32'h10031a74)
`define MLDSA_REG_MLDSA_SIGNATURE_975                                                               (32'h1a74)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_976                                                           (32'h10031a78)
`define MLDSA_REG_MLDSA_SIGNATURE_976                                                               (32'h1a78)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_977                                                           (32'h10031a7c)
`define MLDSA_REG_MLDSA_SIGNATURE_977                                                               (32'h1a7c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_978                                                           (32'h10031a80)
`define MLDSA_REG_MLDSA_SIGNATURE_978                                                               (32'h1a80)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_979                                                           (32'h10031a84)
`define MLDSA_REG_MLDSA_SIGNATURE_979                                                               (32'h1a84)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_980                                                           (32'h10031a88)
`define MLDSA_REG_MLDSA_SIGNATURE_980                                                               (32'h1a88)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_981                                                           (32'h10031a8c)
`define MLDSA_REG_MLDSA_SIGNATURE_981                                                               (32'h1a8c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_982                                                           (32'h10031a90)
`define MLDSA_REG_MLDSA_SIGNATURE_982                                                               (32'h1a90)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_983                                                           (32'h10031a94)
`define MLDSA_REG_MLDSA_SIGNATURE_983                                                               (32'h1a94)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_984                                                           (32'h10031a98)
`define MLDSA_REG_MLDSA_SIGNATURE_984                                                               (32'h1a98)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_985                                                           (32'h10031a9c)
`define MLDSA_REG_MLDSA_SIGNATURE_985                                                               (32'h1a9c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_986                                                           (32'h10031aa0)
`define MLDSA_REG_MLDSA_SIGNATURE_986                                                               (32'h1aa0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_987                                                           (32'h10031aa4)
`define MLDSA_REG_MLDSA_SIGNATURE_987                                                               (32'h1aa4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_988                                                           (32'h10031aa8)
`define MLDSA_REG_MLDSA_SIGNATURE_988                                                               (32'h1aa8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_989                                                           (32'h10031aac)
`define MLDSA_REG_MLDSA_SIGNATURE_989                                                               (32'h1aac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_990                                                           (32'h10031ab0)
`define MLDSA_REG_MLDSA_SIGNATURE_990                                                               (32'h1ab0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_991                                                           (32'h10031ab4)
`define MLDSA_REG_MLDSA_SIGNATURE_991                                                               (32'h1ab4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_992                                                           (32'h10031ab8)
`define MLDSA_REG_MLDSA_SIGNATURE_992                                                               (32'h1ab8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_993                                                           (32'h10031abc)
`define MLDSA_REG_MLDSA_SIGNATURE_993                                                               (32'h1abc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_994                                                           (32'h10031ac0)
`define MLDSA_REG_MLDSA_SIGNATURE_994                                                               (32'h1ac0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_995                                                           (32'h10031ac4)
`define MLDSA_REG_MLDSA_SIGNATURE_995                                                               (32'h1ac4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_996                                                           (32'h10031ac8)
`define MLDSA_REG_MLDSA_SIGNATURE_996                                                               (32'h1ac8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_997                                                           (32'h10031acc)
`define MLDSA_REG_MLDSA_SIGNATURE_997                                                               (32'h1acc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_998                                                           (32'h10031ad0)
`define MLDSA_REG_MLDSA_SIGNATURE_998                                                               (32'h1ad0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_999                                                           (32'h10031ad4)
`define MLDSA_REG_MLDSA_SIGNATURE_999                                                               (32'h1ad4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1000                                                          (32'h10031ad8)
`define MLDSA_REG_MLDSA_SIGNATURE_1000                                                              (32'h1ad8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1001                                                          (32'h10031adc)
`define MLDSA_REG_MLDSA_SIGNATURE_1001                                                              (32'h1adc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1002                                                          (32'h10031ae0)
`define MLDSA_REG_MLDSA_SIGNATURE_1002                                                              (32'h1ae0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1003                                                          (32'h10031ae4)
`define MLDSA_REG_MLDSA_SIGNATURE_1003                                                              (32'h1ae4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1004                                                          (32'h10031ae8)
`define MLDSA_REG_MLDSA_SIGNATURE_1004                                                              (32'h1ae8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1005                                                          (32'h10031aec)
`define MLDSA_REG_MLDSA_SIGNATURE_1005                                                              (32'h1aec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1006                                                          (32'h10031af0)
`define MLDSA_REG_MLDSA_SIGNATURE_1006                                                              (32'h1af0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1007                                                          (32'h10031af4)
`define MLDSA_REG_MLDSA_SIGNATURE_1007                                                              (32'h1af4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1008                                                          (32'h10031af8)
`define MLDSA_REG_MLDSA_SIGNATURE_1008                                                              (32'h1af8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1009                                                          (32'h10031afc)
`define MLDSA_REG_MLDSA_SIGNATURE_1009                                                              (32'h1afc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1010                                                          (32'h10031b00)
`define MLDSA_REG_MLDSA_SIGNATURE_1010                                                              (32'h1b00)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1011                                                          (32'h10031b04)
`define MLDSA_REG_MLDSA_SIGNATURE_1011                                                              (32'h1b04)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1012                                                          (32'h10031b08)
`define MLDSA_REG_MLDSA_SIGNATURE_1012                                                              (32'h1b08)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1013                                                          (32'h10031b0c)
`define MLDSA_REG_MLDSA_SIGNATURE_1013                                                              (32'h1b0c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1014                                                          (32'h10031b10)
`define MLDSA_REG_MLDSA_SIGNATURE_1014                                                              (32'h1b10)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1015                                                          (32'h10031b14)
`define MLDSA_REG_MLDSA_SIGNATURE_1015                                                              (32'h1b14)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1016                                                          (32'h10031b18)
`define MLDSA_REG_MLDSA_SIGNATURE_1016                                                              (32'h1b18)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1017                                                          (32'h10031b1c)
`define MLDSA_REG_MLDSA_SIGNATURE_1017                                                              (32'h1b1c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1018                                                          (32'h10031b20)
`define MLDSA_REG_MLDSA_SIGNATURE_1018                                                              (32'h1b20)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1019                                                          (32'h10031b24)
`define MLDSA_REG_MLDSA_SIGNATURE_1019                                                              (32'h1b24)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1020                                                          (32'h10031b28)
`define MLDSA_REG_MLDSA_SIGNATURE_1020                                                              (32'h1b28)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1021                                                          (32'h10031b2c)
`define MLDSA_REG_MLDSA_SIGNATURE_1021                                                              (32'h1b2c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1022                                                          (32'h10031b30)
`define MLDSA_REG_MLDSA_SIGNATURE_1022                                                              (32'h1b30)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1023                                                          (32'h10031b34)
`define MLDSA_REG_MLDSA_SIGNATURE_1023                                                              (32'h1b34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1024                                                          (32'h10031b38)
`define MLDSA_REG_MLDSA_SIGNATURE_1024                                                              (32'h1b38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1025                                                          (32'h10031b3c)
`define MLDSA_REG_MLDSA_SIGNATURE_1025                                                              (32'h1b3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1026                                                          (32'h10031b40)
`define MLDSA_REG_MLDSA_SIGNATURE_1026                                                              (32'h1b40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1027                                                          (32'h10031b44)
`define MLDSA_REG_MLDSA_SIGNATURE_1027                                                              (32'h1b44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1028                                                          (32'h10031b48)
`define MLDSA_REG_MLDSA_SIGNATURE_1028                                                              (32'h1b48)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1029                                                          (32'h10031b4c)
`define MLDSA_REG_MLDSA_SIGNATURE_1029                                                              (32'h1b4c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1030                                                          (32'h10031b50)
`define MLDSA_REG_MLDSA_SIGNATURE_1030                                                              (32'h1b50)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1031                                                          (32'h10031b54)
`define MLDSA_REG_MLDSA_SIGNATURE_1031                                                              (32'h1b54)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1032                                                          (32'h10031b58)
`define MLDSA_REG_MLDSA_SIGNATURE_1032                                                              (32'h1b58)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1033                                                          (32'h10031b5c)
`define MLDSA_REG_MLDSA_SIGNATURE_1033                                                              (32'h1b5c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1034                                                          (32'h10031b60)
`define MLDSA_REG_MLDSA_SIGNATURE_1034                                                              (32'h1b60)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1035                                                          (32'h10031b64)
`define MLDSA_REG_MLDSA_SIGNATURE_1035                                                              (32'h1b64)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1036                                                          (32'h10031b68)
`define MLDSA_REG_MLDSA_SIGNATURE_1036                                                              (32'h1b68)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1037                                                          (32'h10031b6c)
`define MLDSA_REG_MLDSA_SIGNATURE_1037                                                              (32'h1b6c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1038                                                          (32'h10031b70)
`define MLDSA_REG_MLDSA_SIGNATURE_1038                                                              (32'h1b70)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1039                                                          (32'h10031b74)
`define MLDSA_REG_MLDSA_SIGNATURE_1039                                                              (32'h1b74)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1040                                                          (32'h10031b78)
`define MLDSA_REG_MLDSA_SIGNATURE_1040                                                              (32'h1b78)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1041                                                          (32'h10031b7c)
`define MLDSA_REG_MLDSA_SIGNATURE_1041                                                              (32'h1b7c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1042                                                          (32'h10031b80)
`define MLDSA_REG_MLDSA_SIGNATURE_1042                                                              (32'h1b80)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1043                                                          (32'h10031b84)
`define MLDSA_REG_MLDSA_SIGNATURE_1043                                                              (32'h1b84)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1044                                                          (32'h10031b88)
`define MLDSA_REG_MLDSA_SIGNATURE_1044                                                              (32'h1b88)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1045                                                          (32'h10031b8c)
`define MLDSA_REG_MLDSA_SIGNATURE_1045                                                              (32'h1b8c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1046                                                          (32'h10031b90)
`define MLDSA_REG_MLDSA_SIGNATURE_1046                                                              (32'h1b90)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1047                                                          (32'h10031b94)
`define MLDSA_REG_MLDSA_SIGNATURE_1047                                                              (32'h1b94)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1048                                                          (32'h10031b98)
`define MLDSA_REG_MLDSA_SIGNATURE_1048                                                              (32'h1b98)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1049                                                          (32'h10031b9c)
`define MLDSA_REG_MLDSA_SIGNATURE_1049                                                              (32'h1b9c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1050                                                          (32'h10031ba0)
`define MLDSA_REG_MLDSA_SIGNATURE_1050                                                              (32'h1ba0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1051                                                          (32'h10031ba4)
`define MLDSA_REG_MLDSA_SIGNATURE_1051                                                              (32'h1ba4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1052                                                          (32'h10031ba8)
`define MLDSA_REG_MLDSA_SIGNATURE_1052                                                              (32'h1ba8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1053                                                          (32'h10031bac)
`define MLDSA_REG_MLDSA_SIGNATURE_1053                                                              (32'h1bac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1054                                                          (32'h10031bb0)
`define MLDSA_REG_MLDSA_SIGNATURE_1054                                                              (32'h1bb0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1055                                                          (32'h10031bb4)
`define MLDSA_REG_MLDSA_SIGNATURE_1055                                                              (32'h1bb4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1056                                                          (32'h10031bb8)
`define MLDSA_REG_MLDSA_SIGNATURE_1056                                                              (32'h1bb8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1057                                                          (32'h10031bbc)
`define MLDSA_REG_MLDSA_SIGNATURE_1057                                                              (32'h1bbc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1058                                                          (32'h10031bc0)
`define MLDSA_REG_MLDSA_SIGNATURE_1058                                                              (32'h1bc0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1059                                                          (32'h10031bc4)
`define MLDSA_REG_MLDSA_SIGNATURE_1059                                                              (32'h1bc4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1060                                                          (32'h10031bc8)
`define MLDSA_REG_MLDSA_SIGNATURE_1060                                                              (32'h1bc8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1061                                                          (32'h10031bcc)
`define MLDSA_REG_MLDSA_SIGNATURE_1061                                                              (32'h1bcc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1062                                                          (32'h10031bd0)
`define MLDSA_REG_MLDSA_SIGNATURE_1062                                                              (32'h1bd0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1063                                                          (32'h10031bd4)
`define MLDSA_REG_MLDSA_SIGNATURE_1063                                                              (32'h1bd4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1064                                                          (32'h10031bd8)
`define MLDSA_REG_MLDSA_SIGNATURE_1064                                                              (32'h1bd8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1065                                                          (32'h10031bdc)
`define MLDSA_REG_MLDSA_SIGNATURE_1065                                                              (32'h1bdc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1066                                                          (32'h10031be0)
`define MLDSA_REG_MLDSA_SIGNATURE_1066                                                              (32'h1be0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1067                                                          (32'h10031be4)
`define MLDSA_REG_MLDSA_SIGNATURE_1067                                                              (32'h1be4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1068                                                          (32'h10031be8)
`define MLDSA_REG_MLDSA_SIGNATURE_1068                                                              (32'h1be8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1069                                                          (32'h10031bec)
`define MLDSA_REG_MLDSA_SIGNATURE_1069                                                              (32'h1bec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1070                                                          (32'h10031bf0)
`define MLDSA_REG_MLDSA_SIGNATURE_1070                                                              (32'h1bf0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1071                                                          (32'h10031bf4)
`define MLDSA_REG_MLDSA_SIGNATURE_1071                                                              (32'h1bf4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1072                                                          (32'h10031bf8)
`define MLDSA_REG_MLDSA_SIGNATURE_1072                                                              (32'h1bf8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1073                                                          (32'h10031bfc)
`define MLDSA_REG_MLDSA_SIGNATURE_1073                                                              (32'h1bfc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1074                                                          (32'h10031c00)
`define MLDSA_REG_MLDSA_SIGNATURE_1074                                                              (32'h1c00)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1075                                                          (32'h10031c04)
`define MLDSA_REG_MLDSA_SIGNATURE_1075                                                              (32'h1c04)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1076                                                          (32'h10031c08)
`define MLDSA_REG_MLDSA_SIGNATURE_1076                                                              (32'h1c08)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1077                                                          (32'h10031c0c)
`define MLDSA_REG_MLDSA_SIGNATURE_1077                                                              (32'h1c0c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1078                                                          (32'h10031c10)
`define MLDSA_REG_MLDSA_SIGNATURE_1078                                                              (32'h1c10)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1079                                                          (32'h10031c14)
`define MLDSA_REG_MLDSA_SIGNATURE_1079                                                              (32'h1c14)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1080                                                          (32'h10031c18)
`define MLDSA_REG_MLDSA_SIGNATURE_1080                                                              (32'h1c18)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1081                                                          (32'h10031c1c)
`define MLDSA_REG_MLDSA_SIGNATURE_1081                                                              (32'h1c1c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1082                                                          (32'h10031c20)
`define MLDSA_REG_MLDSA_SIGNATURE_1082                                                              (32'h1c20)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1083                                                          (32'h10031c24)
`define MLDSA_REG_MLDSA_SIGNATURE_1083                                                              (32'h1c24)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1084                                                          (32'h10031c28)
`define MLDSA_REG_MLDSA_SIGNATURE_1084                                                              (32'h1c28)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1085                                                          (32'h10031c2c)
`define MLDSA_REG_MLDSA_SIGNATURE_1085                                                              (32'h1c2c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1086                                                          (32'h10031c30)
`define MLDSA_REG_MLDSA_SIGNATURE_1086                                                              (32'h1c30)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1087                                                          (32'h10031c34)
`define MLDSA_REG_MLDSA_SIGNATURE_1087                                                              (32'h1c34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1088                                                          (32'h10031c38)
`define MLDSA_REG_MLDSA_SIGNATURE_1088                                                              (32'h1c38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1089                                                          (32'h10031c3c)
`define MLDSA_REG_MLDSA_SIGNATURE_1089                                                              (32'h1c3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1090                                                          (32'h10031c40)
`define MLDSA_REG_MLDSA_SIGNATURE_1090                                                              (32'h1c40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1091                                                          (32'h10031c44)
`define MLDSA_REG_MLDSA_SIGNATURE_1091                                                              (32'h1c44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1092                                                          (32'h10031c48)
`define MLDSA_REG_MLDSA_SIGNATURE_1092                                                              (32'h1c48)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1093                                                          (32'h10031c4c)
`define MLDSA_REG_MLDSA_SIGNATURE_1093                                                              (32'h1c4c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1094                                                          (32'h10031c50)
`define MLDSA_REG_MLDSA_SIGNATURE_1094                                                              (32'h1c50)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1095                                                          (32'h10031c54)
`define MLDSA_REG_MLDSA_SIGNATURE_1095                                                              (32'h1c54)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1096                                                          (32'h10031c58)
`define MLDSA_REG_MLDSA_SIGNATURE_1096                                                              (32'h1c58)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1097                                                          (32'h10031c5c)
`define MLDSA_REG_MLDSA_SIGNATURE_1097                                                              (32'h1c5c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1098                                                          (32'h10031c60)
`define MLDSA_REG_MLDSA_SIGNATURE_1098                                                              (32'h1c60)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1099                                                          (32'h10031c64)
`define MLDSA_REG_MLDSA_SIGNATURE_1099                                                              (32'h1c64)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1100                                                          (32'h10031c68)
`define MLDSA_REG_MLDSA_SIGNATURE_1100                                                              (32'h1c68)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1101                                                          (32'h10031c6c)
`define MLDSA_REG_MLDSA_SIGNATURE_1101                                                              (32'h1c6c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1102                                                          (32'h10031c70)
`define MLDSA_REG_MLDSA_SIGNATURE_1102                                                              (32'h1c70)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1103                                                          (32'h10031c74)
`define MLDSA_REG_MLDSA_SIGNATURE_1103                                                              (32'h1c74)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1104                                                          (32'h10031c78)
`define MLDSA_REG_MLDSA_SIGNATURE_1104                                                              (32'h1c78)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1105                                                          (32'h10031c7c)
`define MLDSA_REG_MLDSA_SIGNATURE_1105                                                              (32'h1c7c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1106                                                          (32'h10031c80)
`define MLDSA_REG_MLDSA_SIGNATURE_1106                                                              (32'h1c80)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1107                                                          (32'h10031c84)
`define MLDSA_REG_MLDSA_SIGNATURE_1107                                                              (32'h1c84)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1108                                                          (32'h10031c88)
`define MLDSA_REG_MLDSA_SIGNATURE_1108                                                              (32'h1c88)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1109                                                          (32'h10031c8c)
`define MLDSA_REG_MLDSA_SIGNATURE_1109                                                              (32'h1c8c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1110                                                          (32'h10031c90)
`define MLDSA_REG_MLDSA_SIGNATURE_1110                                                              (32'h1c90)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1111                                                          (32'h10031c94)
`define MLDSA_REG_MLDSA_SIGNATURE_1111                                                              (32'h1c94)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1112                                                          (32'h10031c98)
`define MLDSA_REG_MLDSA_SIGNATURE_1112                                                              (32'h1c98)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1113                                                          (32'h10031c9c)
`define MLDSA_REG_MLDSA_SIGNATURE_1113                                                              (32'h1c9c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1114                                                          (32'h10031ca0)
`define MLDSA_REG_MLDSA_SIGNATURE_1114                                                              (32'h1ca0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1115                                                          (32'h10031ca4)
`define MLDSA_REG_MLDSA_SIGNATURE_1115                                                              (32'h1ca4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1116                                                          (32'h10031ca8)
`define MLDSA_REG_MLDSA_SIGNATURE_1116                                                              (32'h1ca8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1117                                                          (32'h10031cac)
`define MLDSA_REG_MLDSA_SIGNATURE_1117                                                              (32'h1cac)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1118                                                          (32'h10031cb0)
`define MLDSA_REG_MLDSA_SIGNATURE_1118                                                              (32'h1cb0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1119                                                          (32'h10031cb4)
`define MLDSA_REG_MLDSA_SIGNATURE_1119                                                              (32'h1cb4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1120                                                          (32'h10031cb8)
`define MLDSA_REG_MLDSA_SIGNATURE_1120                                                              (32'h1cb8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1121                                                          (32'h10031cbc)
`define MLDSA_REG_MLDSA_SIGNATURE_1121                                                              (32'h1cbc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1122                                                          (32'h10031cc0)
`define MLDSA_REG_MLDSA_SIGNATURE_1122                                                              (32'h1cc0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1123                                                          (32'h10031cc4)
`define MLDSA_REG_MLDSA_SIGNATURE_1123                                                              (32'h1cc4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1124                                                          (32'h10031cc8)
`define MLDSA_REG_MLDSA_SIGNATURE_1124                                                              (32'h1cc8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1125                                                          (32'h10031ccc)
`define MLDSA_REG_MLDSA_SIGNATURE_1125                                                              (32'h1ccc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1126                                                          (32'h10031cd0)
`define MLDSA_REG_MLDSA_SIGNATURE_1126                                                              (32'h1cd0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1127                                                          (32'h10031cd4)
`define MLDSA_REG_MLDSA_SIGNATURE_1127                                                              (32'h1cd4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1128                                                          (32'h10031cd8)
`define MLDSA_REG_MLDSA_SIGNATURE_1128                                                              (32'h1cd8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1129                                                          (32'h10031cdc)
`define MLDSA_REG_MLDSA_SIGNATURE_1129                                                              (32'h1cdc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1130                                                          (32'h10031ce0)
`define MLDSA_REG_MLDSA_SIGNATURE_1130                                                              (32'h1ce0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1131                                                          (32'h10031ce4)
`define MLDSA_REG_MLDSA_SIGNATURE_1131                                                              (32'h1ce4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1132                                                          (32'h10031ce8)
`define MLDSA_REG_MLDSA_SIGNATURE_1132                                                              (32'h1ce8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1133                                                          (32'h10031cec)
`define MLDSA_REG_MLDSA_SIGNATURE_1133                                                              (32'h1cec)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1134                                                          (32'h10031cf0)
`define MLDSA_REG_MLDSA_SIGNATURE_1134                                                              (32'h1cf0)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1135                                                          (32'h10031cf4)
`define MLDSA_REG_MLDSA_SIGNATURE_1135                                                              (32'h1cf4)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1136                                                          (32'h10031cf8)
`define MLDSA_REG_MLDSA_SIGNATURE_1136                                                              (32'h1cf8)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1137                                                          (32'h10031cfc)
`define MLDSA_REG_MLDSA_SIGNATURE_1137                                                              (32'h1cfc)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1138                                                          (32'h10031d00)
`define MLDSA_REG_MLDSA_SIGNATURE_1138                                                              (32'h1d00)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1139                                                          (32'h10031d04)
`define MLDSA_REG_MLDSA_SIGNATURE_1139                                                              (32'h1d04)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1140                                                          (32'h10031d08)
`define MLDSA_REG_MLDSA_SIGNATURE_1140                                                              (32'h1d08)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1141                                                          (32'h10031d0c)
`define MLDSA_REG_MLDSA_SIGNATURE_1141                                                              (32'h1d0c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1142                                                          (32'h10031d10)
`define MLDSA_REG_MLDSA_SIGNATURE_1142                                                              (32'h1d10)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1143                                                          (32'h10031d14)
`define MLDSA_REG_MLDSA_SIGNATURE_1143                                                              (32'h1d14)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1144                                                          (32'h10031d18)
`define MLDSA_REG_MLDSA_SIGNATURE_1144                                                              (32'h1d18)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1145                                                          (32'h10031d1c)
`define MLDSA_REG_MLDSA_SIGNATURE_1145                                                              (32'h1d1c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1146                                                          (32'h10031d20)
`define MLDSA_REG_MLDSA_SIGNATURE_1146                                                              (32'h1d20)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1147                                                          (32'h10031d24)
`define MLDSA_REG_MLDSA_SIGNATURE_1147                                                              (32'h1d24)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1148                                                          (32'h10031d28)
`define MLDSA_REG_MLDSA_SIGNATURE_1148                                                              (32'h1d28)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1149                                                          (32'h10031d2c)
`define MLDSA_REG_MLDSA_SIGNATURE_1149                                                              (32'h1d2c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1150                                                          (32'h10031d30)
`define MLDSA_REG_MLDSA_SIGNATURE_1150                                                              (32'h1d30)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1151                                                          (32'h10031d34)
`define MLDSA_REG_MLDSA_SIGNATURE_1151                                                              (32'h1d34)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1152                                                          (32'h10031d38)
`define MLDSA_REG_MLDSA_SIGNATURE_1152                                                              (32'h1d38)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1153                                                          (32'h10031d3c)
`define MLDSA_REG_MLDSA_SIGNATURE_1153                                                              (32'h1d3c)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1154                                                          (32'h10031d40)
`define MLDSA_REG_MLDSA_SIGNATURE_1154                                                              (32'h1d40)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1155                                                          (32'h10031d44)
`define MLDSA_REG_MLDSA_SIGNATURE_1155                                                              (32'h1d44)
`define CLP_MLDSA_REG_MLDSA_SIGNATURE_1156                                                          (32'h10031d48)
`define MLDSA_REG_MLDSA_SIGNATURE_1156                                                              (32'h1d48)
`define CLP_MLDSA_REG_MLDSA_PRIVKEY_OUT_BASE_ADDR                                                   (32'h10032000)
`define CLP_MLDSA_REG_MLDSA_PRIVKEY_OUT_END_ADDR                                                    (32'h1003331f)
`define CLP_MLDSA_REG_MLDSA_PRIVKEY_IN_BASE_ADDR                                                    (32'h10034000)
`define CLP_MLDSA_REG_MLDSA_PRIVKEY_IN_END_ADDR                                                     (32'h1003531f)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_START                                                           (32'h10036000)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                (32'h10036000)
`define MLDSA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                    (32'h6000)
`define MLDSA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                       (0)
`define MLDSA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                      (32'h1)
`define MLDSA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                       (1)
`define MLDSA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                      (32'h2)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                 (32'h10036004)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                     (32'h6004)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_LOW                               (0)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_MASK                              (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                 (32'h10036008)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                     (32'h6008)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                               (0)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                              (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                             (32'h1003600c)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                 (32'h600c)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                     (0)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                    (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                             (32'h10036010)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                 (32'h6010)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                     (0)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                    (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                           (32'h10036014)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                               (32'h6014)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_LOW                        (0)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_MASK                       (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                           (32'h10036018)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                               (32'h6018)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                        (0)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                       (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                               (32'h1003601c)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                   (32'h601c)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_LOW                           (0)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_MASK                          (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                               (32'h10036020)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                   (32'h6020)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                           (0)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                          (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                     (32'h10036100)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                         (32'h6100)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                     (32'h10036180)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                         (32'h6180)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                (32'h10036200)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                    (32'h6200)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_LOW                          (0)
`define MLDSA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_MASK                         (32'h1)
`define CLP_MLDSA_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                (32'h10036204)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                    (32'h6204)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                          (0)
`define MLDSA_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                         (32'h1)
`define CLP_SPI_HOST_REG_BASE_ADDR                                                                  (32'h20000000)
`define CLP_SPI_HOST_REG_INTERRUPT_STATE                                                            (32'h20000000)
`define SPI_HOST_REG_INTERRUPT_STATE                                                                (32'h0)
`define SPI_HOST_REG_INTERRUPT_STATE_ERROR_LOW                                                      (0)
`define SPI_HOST_REG_INTERRUPT_STATE_ERROR_MASK                                                     (32'h1)
`define SPI_HOST_REG_INTERRUPT_STATE_SPI_EVENT_LOW                                                  (1)
`define SPI_HOST_REG_INTERRUPT_STATE_SPI_EVENT_MASK                                                 (32'h2)
`define CLP_SPI_HOST_REG_INTERRUPT_ENABLE                                                           (32'h20000004)
`define SPI_HOST_REG_INTERRUPT_ENABLE                                                               (32'h4)
`define SPI_HOST_REG_INTERRUPT_ENABLE_ERROR_LOW                                                     (0)
`define SPI_HOST_REG_INTERRUPT_ENABLE_ERROR_MASK                                                    (32'h1)
`define SPI_HOST_REG_INTERRUPT_ENABLE_SPI_EVENT_LOW                                                 (1)
`define SPI_HOST_REG_INTERRUPT_ENABLE_SPI_EVENT_MASK                                                (32'h2)
`define CLP_SPI_HOST_REG_INTERRUPT_TEST                                                             (32'h20000008)
`define SPI_HOST_REG_INTERRUPT_TEST                                                                 (32'h8)
`define SPI_HOST_REG_INTERRUPT_TEST_ERROR_LOW                                                       (0)
`define SPI_HOST_REG_INTERRUPT_TEST_ERROR_MASK                                                      (32'h1)
`define SPI_HOST_REG_INTERRUPT_TEST_SPI_EVENT_LOW                                                   (1)
`define SPI_HOST_REG_INTERRUPT_TEST_SPI_EVENT_MASK                                                  (32'h2)
`define CLP_SPI_HOST_REG_ALERT_TEST                                                                 (32'h2000000c)
`define SPI_HOST_REG_ALERT_TEST                                                                     (32'hc)
`define SPI_HOST_REG_ALERT_TEST_FATAL_FAULT_LOW                                                     (0)
`define SPI_HOST_REG_ALERT_TEST_FATAL_FAULT_MASK                                                    (32'h1)
`define CLP_SPI_HOST_REG_CONTROL                                                                    (32'h20000010)
`define SPI_HOST_REG_CONTROL                                                                        (32'h10)
`define SPI_HOST_REG_CONTROL_RX_WATERMARK_LOW                                                       (0)
`define SPI_HOST_REG_CONTROL_RX_WATERMARK_MASK                                                      (32'hff)
`define SPI_HOST_REG_CONTROL_TX_WATERMARK_LOW                                                       (8)
`define SPI_HOST_REG_CONTROL_TX_WATERMARK_MASK                                                      (32'hff00)
`define SPI_HOST_REG_CONTROL_OUTPUT_EN_LOW                                                          (29)
`define SPI_HOST_REG_CONTROL_OUTPUT_EN_MASK                                                         (32'h20000000)
`define SPI_HOST_REG_CONTROL_SW_RST_LOW                                                             (30)
`define SPI_HOST_REG_CONTROL_SW_RST_MASK                                                            (32'h40000000)
`define SPI_HOST_REG_CONTROL_SPIEN_LOW                                                              (31)
`define SPI_HOST_REG_CONTROL_SPIEN_MASK                                                             (32'h80000000)
`define CLP_SPI_HOST_REG_STATUS                                                                     (32'h20000014)
`define SPI_HOST_REG_STATUS                                                                         (32'h14)
`define SPI_HOST_REG_STATUS_TXQD_LOW                                                                (0)
`define SPI_HOST_REG_STATUS_TXQD_MASK                                                               (32'hff)
`define SPI_HOST_REG_STATUS_RXQD_LOW                                                                (8)
`define SPI_HOST_REG_STATUS_RXQD_MASK                                                               (32'hff00)
`define SPI_HOST_REG_STATUS_CMDQD_LOW                                                               (16)
`define SPI_HOST_REG_STATUS_CMDQD_MASK                                                              (32'hf0000)
`define SPI_HOST_REG_STATUS_RXWM_LOW                                                                (20)
`define SPI_HOST_REG_STATUS_RXWM_MASK                                                               (32'h100000)
`define SPI_HOST_REG_STATUS_BYTEORDER_LOW                                                           (22)
`define SPI_HOST_REG_STATUS_BYTEORDER_MASK                                                          (32'h400000)
`define SPI_HOST_REG_STATUS_RXSTALL_LOW                                                             (23)
`define SPI_HOST_REG_STATUS_RXSTALL_MASK                                                            (32'h800000)
`define SPI_HOST_REG_STATUS_RXEMPTY_LOW                                                             (24)
`define SPI_HOST_REG_STATUS_RXEMPTY_MASK                                                            (32'h1000000)
`define SPI_HOST_REG_STATUS_RXFULL_LOW                                                              (25)
`define SPI_HOST_REG_STATUS_RXFULL_MASK                                                             (32'h2000000)
`define SPI_HOST_REG_STATUS_TXWM_LOW                                                                (26)
`define SPI_HOST_REG_STATUS_TXWM_MASK                                                               (32'h4000000)
`define SPI_HOST_REG_STATUS_TXSTALL_LOW                                                             (27)
`define SPI_HOST_REG_STATUS_TXSTALL_MASK                                                            (32'h8000000)
`define SPI_HOST_REG_STATUS_TXEMPTY_LOW                                                             (28)
`define SPI_HOST_REG_STATUS_TXEMPTY_MASK                                                            (32'h10000000)
`define SPI_HOST_REG_STATUS_TXFULL_LOW                                                              (29)
`define SPI_HOST_REG_STATUS_TXFULL_MASK                                                             (32'h20000000)
`define SPI_HOST_REG_STATUS_ACTIVE_LOW                                                              (30)
`define SPI_HOST_REG_STATUS_ACTIVE_MASK                                                             (32'h40000000)
`define SPI_HOST_REG_STATUS_READY_LOW                                                               (31)
`define SPI_HOST_REG_STATUS_READY_MASK                                                              (32'h80000000)
`define CLP_SPI_HOST_REG_CONFIGOPTS_0                                                               (32'h20000018)
`define SPI_HOST_REG_CONFIGOPTS_0                                                                   (32'h18)
`define SPI_HOST_REG_CONFIGOPTS_0_CLKDIV_LOW                                                        (0)
`define SPI_HOST_REG_CONFIGOPTS_0_CLKDIV_MASK                                                       (32'hffff)
`define SPI_HOST_REG_CONFIGOPTS_0_CSNIDLE_LOW                                                       (16)
`define SPI_HOST_REG_CONFIGOPTS_0_CSNIDLE_MASK                                                      (32'hf0000)
`define SPI_HOST_REG_CONFIGOPTS_0_CSNTRAIL_LOW                                                      (20)
`define SPI_HOST_REG_CONFIGOPTS_0_CSNTRAIL_MASK                                                     (32'hf00000)
`define SPI_HOST_REG_CONFIGOPTS_0_CSNLEAD_LOW                                                       (24)
`define SPI_HOST_REG_CONFIGOPTS_0_CSNLEAD_MASK                                                      (32'hf000000)
`define SPI_HOST_REG_CONFIGOPTS_0_FULLCYC_LOW                                                       (29)
`define SPI_HOST_REG_CONFIGOPTS_0_FULLCYC_MASK                                                      (32'h20000000)
`define SPI_HOST_REG_CONFIGOPTS_0_CPHA_LOW                                                          (30)
`define SPI_HOST_REG_CONFIGOPTS_0_CPHA_MASK                                                         (32'h40000000)
`define SPI_HOST_REG_CONFIGOPTS_0_CPOL_LOW                                                          (31)
`define SPI_HOST_REG_CONFIGOPTS_0_CPOL_MASK                                                         (32'h80000000)
`define CLP_SPI_HOST_REG_CONFIGOPTS_1                                                               (32'h2000001c)
`define SPI_HOST_REG_CONFIGOPTS_1                                                                   (32'h1c)
`define SPI_HOST_REG_CONFIGOPTS_1_CLKDIV_LOW                                                        (0)
`define SPI_HOST_REG_CONFIGOPTS_1_CLKDIV_MASK                                                       (32'hffff)
`define SPI_HOST_REG_CONFIGOPTS_1_CSNIDLE_LOW                                                       (16)
`define SPI_HOST_REG_CONFIGOPTS_1_CSNIDLE_MASK                                                      (32'hf0000)
`define SPI_HOST_REG_CONFIGOPTS_1_CSNTRAIL_LOW                                                      (20)
`define SPI_HOST_REG_CONFIGOPTS_1_CSNTRAIL_MASK                                                     (32'hf00000)
`define SPI_HOST_REG_CONFIGOPTS_1_CSNLEAD_LOW                                                       (24)
`define SPI_HOST_REG_CONFIGOPTS_1_CSNLEAD_MASK                                                      (32'hf000000)
`define SPI_HOST_REG_CONFIGOPTS_1_FULLCYC_LOW                                                       (29)
`define SPI_HOST_REG_CONFIGOPTS_1_FULLCYC_MASK                                                      (32'h20000000)
`define SPI_HOST_REG_CONFIGOPTS_1_CPHA_LOW                                                          (30)
`define SPI_HOST_REG_CONFIGOPTS_1_CPHA_MASK                                                         (32'h40000000)
`define SPI_HOST_REG_CONFIGOPTS_1_CPOL_LOW                                                          (31)
`define SPI_HOST_REG_CONFIGOPTS_1_CPOL_MASK                                                         (32'h80000000)
`define CLP_SPI_HOST_REG_CSID                                                                       (32'h20000020)
`define SPI_HOST_REG_CSID                                                                           (32'h20)
`define CLP_SPI_HOST_REG_COMMAND                                                                    (32'h20000024)
`define SPI_HOST_REG_COMMAND                                                                        (32'h24)
`define SPI_HOST_REG_COMMAND_LEN_LOW                                                                (0)
`define SPI_HOST_REG_COMMAND_LEN_MASK                                                               (32'h1ff)
`define SPI_HOST_REG_COMMAND_CSAAT_LOW                                                              (9)
`define SPI_HOST_REG_COMMAND_CSAAT_MASK                                                             (32'h200)
`define SPI_HOST_REG_COMMAND_SPEED_LOW                                                              (10)
`define SPI_HOST_REG_COMMAND_SPEED_MASK                                                             (32'hc00)
`define SPI_HOST_REG_COMMAND_DIRECTION_LOW                                                          (12)
`define SPI_HOST_REG_COMMAND_DIRECTION_MASK                                                         (32'h3000)
`define CLP_SPI_HOST_REG_RXDATA                                                                     (32'h20000028)
`define SPI_HOST_REG_RXDATA                                                                         (32'h28)
`define CLP_SPI_HOST_REG_TXDATA                                                                     (32'h2000002c)
`define SPI_HOST_REG_TXDATA                                                                         (32'h2c)
`define CLP_SPI_HOST_REG_ERROR_ENABLE                                                               (32'h20000030)
`define SPI_HOST_REG_ERROR_ENABLE                                                                   (32'h30)
`define SPI_HOST_REG_ERROR_ENABLE_CMDBUSY_LOW                                                       (0)
`define SPI_HOST_REG_ERROR_ENABLE_CMDBUSY_MASK                                                      (32'h1)
`define SPI_HOST_REG_ERROR_ENABLE_OVERFLOW_LOW                                                      (1)
`define SPI_HOST_REG_ERROR_ENABLE_OVERFLOW_MASK                                                     (32'h2)
`define SPI_HOST_REG_ERROR_ENABLE_UNDERFLOW_LOW                                                     (2)
`define SPI_HOST_REG_ERROR_ENABLE_UNDERFLOW_MASK                                                    (32'h4)
`define SPI_HOST_REG_ERROR_ENABLE_CMDINVAL_LOW                                                      (3)
`define SPI_HOST_REG_ERROR_ENABLE_CMDINVAL_MASK                                                     (32'h8)
`define SPI_HOST_REG_ERROR_ENABLE_CSIDINVAL_LOW                                                     (4)
`define SPI_HOST_REG_ERROR_ENABLE_CSIDINVAL_MASK                                                    (32'h10)
`define CLP_SPI_HOST_REG_ERROR_STATUS                                                               (32'h20000034)
`define SPI_HOST_REG_ERROR_STATUS                                                                   (32'h34)
`define SPI_HOST_REG_ERROR_STATUS_CMDBUSY_LOW                                                       (0)
`define SPI_HOST_REG_ERROR_STATUS_CMDBUSY_MASK                                                      (32'h1)
`define SPI_HOST_REG_ERROR_STATUS_OVERFLOW_LOW                                                      (1)
`define SPI_HOST_REG_ERROR_STATUS_OVERFLOW_MASK                                                     (32'h2)
`define SPI_HOST_REG_ERROR_STATUS_UNDERFLOW_LOW                                                     (2)
`define SPI_HOST_REG_ERROR_STATUS_UNDERFLOW_MASK                                                    (32'h4)
`define SPI_HOST_REG_ERROR_STATUS_CMDINVAL_LOW                                                      (3)
`define SPI_HOST_REG_ERROR_STATUS_CMDINVAL_MASK                                                     (32'h8)
`define SPI_HOST_REG_ERROR_STATUS_CSIDINVAL_LOW                                                     (4)
`define SPI_HOST_REG_ERROR_STATUS_CSIDINVAL_MASK                                                    (32'h10)
`define SPI_HOST_REG_ERROR_STATUS_ACCESSINVAL_LOW                                                   (5)
`define SPI_HOST_REG_ERROR_STATUS_ACCESSINVAL_MASK                                                  (32'h20)
`define CLP_SPI_HOST_REG_EVENT_ENABLE                                                               (32'h20000038)
`define SPI_HOST_REG_EVENT_ENABLE                                                                   (32'h38)
`define SPI_HOST_REG_EVENT_ENABLE_RXFULL_LOW                                                        (0)
`define SPI_HOST_REG_EVENT_ENABLE_RXFULL_MASK                                                       (32'h1)
`define SPI_HOST_REG_EVENT_ENABLE_TXEMPTY_LOW                                                       (1)
`define SPI_HOST_REG_EVENT_ENABLE_TXEMPTY_MASK                                                      (32'h2)
`define SPI_HOST_REG_EVENT_ENABLE_RXWM_LOW                                                          (2)
`define SPI_HOST_REG_EVENT_ENABLE_RXWM_MASK                                                         (32'h4)
`define SPI_HOST_REG_EVENT_ENABLE_TXWM_LOW                                                          (3)
`define SPI_HOST_REG_EVENT_ENABLE_TXWM_MASK                                                         (32'h8)
`define SPI_HOST_REG_EVENT_ENABLE_READY_LOW                                                         (4)
`define SPI_HOST_REG_EVENT_ENABLE_READY_MASK                                                        (32'h10)
`define SPI_HOST_REG_EVENT_ENABLE_IDLE_LOW                                                          (5)
`define SPI_HOST_REG_EVENT_ENABLE_IDLE_MASK                                                         (32'h20)
`define CLP_UART_BASE_ADDR                                                                          (32'h20001000)
`define CLP_UART_INTERRUPT_STATE                                                                    (32'h20001000)
`define UART_INTERRUPT_STATE                                                                        (32'h0)
`define UART_INTERRUPT_STATE_TX_WATERMARK_LOW                                                       (0)
`define UART_INTERRUPT_STATE_TX_WATERMARK_MASK                                                      (32'h1)
`define UART_INTERRUPT_STATE_RX_WATERMARK_LOW                                                       (1)
`define UART_INTERRUPT_STATE_RX_WATERMARK_MASK                                                      (32'h2)
`define UART_INTERRUPT_STATE_TX_EMPTY_LOW                                                           (2)
`define UART_INTERRUPT_STATE_TX_EMPTY_MASK                                                          (32'h4)
`define UART_INTERRUPT_STATE_RX_OVERFLOW_LOW                                                        (3)
`define UART_INTERRUPT_STATE_RX_OVERFLOW_MASK                                                       (32'h8)
`define UART_INTERRUPT_STATE_RX_FRAME_ERR_LOW                                                       (4)
`define UART_INTERRUPT_STATE_RX_FRAME_ERR_MASK                                                      (32'h10)
`define UART_INTERRUPT_STATE_RX_BREAK_ERR_LOW                                                       (5)
`define UART_INTERRUPT_STATE_RX_BREAK_ERR_MASK                                                      (32'h20)
`define UART_INTERRUPT_STATE_RX_TIMEOUT_LOW                                                         (6)
`define UART_INTERRUPT_STATE_RX_TIMEOUT_MASK                                                        (32'h40)
`define UART_INTERRUPT_STATE_RX_PARITY_ERR_LOW                                                      (7)
`define UART_INTERRUPT_STATE_RX_PARITY_ERR_MASK                                                     (32'h80)
`define CLP_UART_INTERRUPT_ENABLE                                                                   (32'h20001004)
`define UART_INTERRUPT_ENABLE                                                                       (32'h4)
`define UART_INTERRUPT_ENABLE_TX_WATERMARK_LOW                                                      (0)
`define UART_INTERRUPT_ENABLE_TX_WATERMARK_MASK                                                     (32'h1)
`define UART_INTERRUPT_ENABLE_RX_WATERMARK_LOW                                                      (1)
`define UART_INTERRUPT_ENABLE_RX_WATERMARK_MASK                                                     (32'h2)
`define UART_INTERRUPT_ENABLE_TX_EMPTY_LOW                                                          (2)
`define UART_INTERRUPT_ENABLE_TX_EMPTY_MASK                                                         (32'h4)
`define UART_INTERRUPT_ENABLE_RX_OVERFLOW_LOW                                                       (3)
`define UART_INTERRUPT_ENABLE_RX_OVERFLOW_MASK                                                      (32'h8)
`define UART_INTERRUPT_ENABLE_RX_FRAME_ERR_LOW                                                      (4)
`define UART_INTERRUPT_ENABLE_RX_FRAME_ERR_MASK                                                     (32'h10)
`define UART_INTERRUPT_ENABLE_RX_BREAK_ERR_LOW                                                      (5)
`define UART_INTERRUPT_ENABLE_RX_BREAK_ERR_MASK                                                     (32'h20)
`define UART_INTERRUPT_ENABLE_RX_TIMEOUT_LOW                                                        (6)
`define UART_INTERRUPT_ENABLE_RX_TIMEOUT_MASK                                                       (32'h40)
`define UART_INTERRUPT_ENABLE_RX_PARITY_ERR_LOW                                                     (7)
`define UART_INTERRUPT_ENABLE_RX_PARITY_ERR_MASK                                                    (32'h80)
`define CLP_UART_INTERRUPT_TEST                                                                     (32'h20001008)
`define UART_INTERRUPT_TEST                                                                         (32'h8)
`define UART_INTERRUPT_TEST_TX_WATERMARK_LOW                                                        (0)
`define UART_INTERRUPT_TEST_TX_WATERMARK_MASK                                                       (32'h1)
`define UART_INTERRUPT_TEST_RX_WATERMARK_LOW                                                        (1)
`define UART_INTERRUPT_TEST_RX_WATERMARK_MASK                                                       (32'h2)
`define UART_INTERRUPT_TEST_TX_EMPTY_LOW                                                            (2)
`define UART_INTERRUPT_TEST_TX_EMPTY_MASK                                                           (32'h4)
`define UART_INTERRUPT_TEST_RX_OVERFLOW_LOW                                                         (3)
`define UART_INTERRUPT_TEST_RX_OVERFLOW_MASK                                                        (32'h8)
`define UART_INTERRUPT_TEST_RX_FRAME_ERR_LOW                                                        (4)
`define UART_INTERRUPT_TEST_RX_FRAME_ERR_MASK                                                       (32'h10)
`define UART_INTERRUPT_TEST_RX_BREAK_ERR_LOW                                                        (5)
`define UART_INTERRUPT_TEST_RX_BREAK_ERR_MASK                                                       (32'h20)
`define UART_INTERRUPT_TEST_RX_TIMEOUT_LOW                                                          (6)
`define UART_INTERRUPT_TEST_RX_TIMEOUT_MASK                                                         (32'h40)
`define UART_INTERRUPT_TEST_RX_PARITY_ERR_LOW                                                       (7)
`define UART_INTERRUPT_TEST_RX_PARITY_ERR_MASK                                                      (32'h80)
`define CLP_UART_ALERT_TEST                                                                         (32'h2000100c)
`define UART_ALERT_TEST                                                                             (32'hc)
`define UART_ALERT_TEST_FATAL_FAULT_LOW                                                             (0)
`define UART_ALERT_TEST_FATAL_FAULT_MASK                                                            (32'h1)
`define CLP_UART_CTRL                                                                               (32'h20001010)
`define UART_CTRL                                                                                   (32'h10)
`define UART_CTRL_TX_LOW                                                                            (0)
`define UART_CTRL_TX_MASK                                                                           (32'h1)
`define UART_CTRL_RX_LOW                                                                            (1)
`define UART_CTRL_RX_MASK                                                                           (32'h2)
`define UART_CTRL_NF_LOW                                                                            (2)
`define UART_CTRL_NF_MASK                                                                           (32'h4)
`define UART_CTRL_SLPBK_LOW                                                                         (4)
`define UART_CTRL_SLPBK_MASK                                                                        (32'h10)
`define UART_CTRL_LLPBK_LOW                                                                         (5)
`define UART_CTRL_LLPBK_MASK                                                                        (32'h20)
`define UART_CTRL_PARITY_EN_LOW                                                                     (6)
`define UART_CTRL_PARITY_EN_MASK                                                                    (32'h40)
`define UART_CTRL_PARITY_ODD_LOW                                                                    (7)
`define UART_CTRL_PARITY_ODD_MASK                                                                   (32'h80)
`define UART_CTRL_RXBLVL_LOW                                                                        (8)
`define UART_CTRL_RXBLVL_MASK                                                                       (32'h300)
`define UART_CTRL_NCO_LOW                                                                           (16)
`define UART_CTRL_NCO_MASK                                                                          (32'hffff0000)
`define CLP_UART_STATUS                                                                             (32'h20001014)
`define UART_STATUS                                                                                 (32'h14)
`define UART_STATUS_TXFULL_LOW                                                                      (0)
`define UART_STATUS_TXFULL_MASK                                                                     (32'h1)
`define UART_STATUS_RXFULL_LOW                                                                      (1)
`define UART_STATUS_RXFULL_MASK                                                                     (32'h2)
`define UART_STATUS_TXEMPTY_LOW                                                                     (2)
`define UART_STATUS_TXEMPTY_MASK                                                                    (32'h4)
`define UART_STATUS_TXIDLE_LOW                                                                      (3)
`define UART_STATUS_TXIDLE_MASK                                                                     (32'h8)
`define UART_STATUS_RXIDLE_LOW                                                                      (4)
`define UART_STATUS_RXIDLE_MASK                                                                     (32'h10)
`define UART_STATUS_RXEMPTY_LOW                                                                     (5)
`define UART_STATUS_RXEMPTY_MASK                                                                    (32'h20)
`define CLP_UART_RDATA                                                                              (32'h20001018)
`define UART_RDATA                                                                                  (32'h18)
`define UART_RDATA_RDATA_LOW                                                                        (0)
`define UART_RDATA_RDATA_MASK                                                                       (32'hff)
`define CLP_UART_WDATA                                                                              (32'h2000101c)
`define UART_WDATA                                                                                  (32'h1c)
`define UART_WDATA_WDATA_LOW                                                                        (0)
`define UART_WDATA_WDATA_MASK                                                                       (32'hff)
`define CLP_UART_FIFO_CTRL                                                                          (32'h20001020)
`define UART_FIFO_CTRL                                                                              (32'h20)
`define UART_FIFO_CTRL_RXRST_LOW                                                                    (0)
`define UART_FIFO_CTRL_RXRST_MASK                                                                   (32'h1)
`define UART_FIFO_CTRL_TXRST_LOW                                                                    (1)
`define UART_FIFO_CTRL_TXRST_MASK                                                                   (32'h2)
`define UART_FIFO_CTRL_RXILVL_LOW                                                                   (2)
`define UART_FIFO_CTRL_RXILVL_MASK                                                                  (32'h1c)
`define UART_FIFO_CTRL_TXILVL_LOW                                                                   (5)
`define UART_FIFO_CTRL_TXILVL_MASK                                                                  (32'h60)
`define CLP_UART_FIFO_STATUS                                                                        (32'h20001024)
`define UART_FIFO_STATUS                                                                            (32'h24)
`define UART_FIFO_STATUS_TXLVL_LOW                                                                  (0)
`define UART_FIFO_STATUS_TXLVL_MASK                                                                 (32'h3f)
`define UART_FIFO_STATUS_RXLVL_LOW                                                                  (16)
`define UART_FIFO_STATUS_RXLVL_MASK                                                                 (32'h3f0000)
`define CLP_UART_OVRD                                                                               (32'h20001028)
`define UART_OVRD                                                                                   (32'h28)
`define UART_OVRD_TXEN_LOW                                                                          (0)
`define UART_OVRD_TXEN_MASK                                                                         (32'h1)
`define UART_OVRD_TXVAL_LOW                                                                         (1)
`define UART_OVRD_TXVAL_MASK                                                                        (32'h2)
`define CLP_UART_VAL                                                                                (32'h2000102c)
`define UART_VAL                                                                                    (32'h2c)
`define UART_VAL_RX_LOW                                                                             (0)
`define UART_VAL_RX_MASK                                                                            (32'hffff)
`define CLP_UART_TIMEOUT_CTRL                                                                       (32'h20001030)
`define UART_TIMEOUT_CTRL                                                                           (32'h30)
`define UART_TIMEOUT_CTRL_VAL_LOW                                                                   (0)
`define UART_TIMEOUT_CTRL_VAL_MASK                                                                  (32'hffffff)
`define UART_TIMEOUT_CTRL_EN_LOW                                                                    (31)
`define UART_TIMEOUT_CTRL_EN_MASK                                                                   (32'h80000000)
`define CLP_CSRNG_REG_BASE_ADDR                                                                     (32'h20002000)
`define CLP_CSRNG_REG_INTERRUPT_STATE                                                               (32'h20002000)
`define CSRNG_REG_INTERRUPT_STATE                                                                   (32'h0)
`define CSRNG_REG_INTERRUPT_STATE_CS_CMD_REQ_DONE_LOW                                               (0)
`define CSRNG_REG_INTERRUPT_STATE_CS_CMD_REQ_DONE_MASK                                              (32'h1)
`define CSRNG_REG_INTERRUPT_STATE_CS_ENTROPY_REQ_LOW                                                (1)
`define CSRNG_REG_INTERRUPT_STATE_CS_ENTROPY_REQ_MASK                                               (32'h2)
`define CSRNG_REG_INTERRUPT_STATE_CS_HW_INST_EXC_LOW                                                (2)
`define CSRNG_REG_INTERRUPT_STATE_CS_HW_INST_EXC_MASK                                               (32'h4)
`define CSRNG_REG_INTERRUPT_STATE_CS_FATAL_ERR_LOW                                                  (3)
`define CSRNG_REG_INTERRUPT_STATE_CS_FATAL_ERR_MASK                                                 (32'h8)
`define CLP_CSRNG_REG_INTERRUPT_ENABLE                                                              (32'h20002004)
`define CSRNG_REG_INTERRUPT_ENABLE                                                                  (32'h4)
`define CSRNG_REG_INTERRUPT_ENABLE_CS_CMD_REQ_DONE_LOW                                              (0)
`define CSRNG_REG_INTERRUPT_ENABLE_CS_CMD_REQ_DONE_MASK                                             (32'h1)
`define CSRNG_REG_INTERRUPT_ENABLE_CS_ENTROPY_REQ_LOW                                               (1)
`define CSRNG_REG_INTERRUPT_ENABLE_CS_ENTROPY_REQ_MASK                                              (32'h2)
`define CSRNG_REG_INTERRUPT_ENABLE_CS_HW_INST_EXC_LOW                                               (2)
`define CSRNG_REG_INTERRUPT_ENABLE_CS_HW_INST_EXC_MASK                                              (32'h4)
`define CSRNG_REG_INTERRUPT_ENABLE_CS_FATAL_ERR_LOW                                                 (3)
`define CSRNG_REG_INTERRUPT_ENABLE_CS_FATAL_ERR_MASK                                                (32'h8)
`define CLP_CSRNG_REG_INTERRUPT_TEST                                                                (32'h20002008)
`define CSRNG_REG_INTERRUPT_TEST                                                                    (32'h8)
`define CSRNG_REG_INTERRUPT_TEST_CS_CMD_REQ_DONE_LOW                                                (0)
`define CSRNG_REG_INTERRUPT_TEST_CS_CMD_REQ_DONE_MASK                                               (32'h1)
`define CSRNG_REG_INTERRUPT_TEST_CS_ENTROPY_REQ_LOW                                                 (1)
`define CSRNG_REG_INTERRUPT_TEST_CS_ENTROPY_REQ_MASK                                                (32'h2)
`define CSRNG_REG_INTERRUPT_TEST_CS_HW_INST_EXC_LOW                                                 (2)
`define CSRNG_REG_INTERRUPT_TEST_CS_HW_INST_EXC_MASK                                                (32'h4)
`define CSRNG_REG_INTERRUPT_TEST_CS_FATAL_ERR_LOW                                                   (3)
`define CSRNG_REG_INTERRUPT_TEST_CS_FATAL_ERR_MASK                                                  (32'h8)
`define CLP_CSRNG_REG_ALERT_TEST                                                                    (32'h2000200c)
`define CSRNG_REG_ALERT_TEST                                                                        (32'hc)
`define CSRNG_REG_ALERT_TEST_RECOV_ALERT_LOW                                                        (0)
`define CSRNG_REG_ALERT_TEST_RECOV_ALERT_MASK                                                       (32'h1)
`define CSRNG_REG_ALERT_TEST_FATAL_ALERT_LOW                                                        (1)
`define CSRNG_REG_ALERT_TEST_FATAL_ALERT_MASK                                                       (32'h2)
`define CLP_CSRNG_REG_REGWEN                                                                        (32'h20002010)
`define CSRNG_REG_REGWEN                                                                            (32'h10)
`define CSRNG_REG_REGWEN_REGWEN_LOW                                                                 (0)
`define CSRNG_REG_REGWEN_REGWEN_MASK                                                                (32'h1)
`define CLP_CSRNG_REG_CTRL                                                                          (32'h20002014)
`define CSRNG_REG_CTRL                                                                              (32'h14)
`define CSRNG_REG_CTRL_ENABLE_LOW                                                                   (0)
`define CSRNG_REG_CTRL_ENABLE_MASK                                                                  (32'hf)
`define CSRNG_REG_CTRL_SW_APP_ENABLE_LOW                                                            (4)
`define CSRNG_REG_CTRL_SW_APP_ENABLE_MASK                                                           (32'hf0)
`define CSRNG_REG_CTRL_READ_INT_STATE_LOW                                                           (8)
`define CSRNG_REG_CTRL_READ_INT_STATE_MASK                                                          (32'hf00)
`define CLP_CSRNG_REG_CMD_REQ                                                                       (32'h20002018)
`define CSRNG_REG_CMD_REQ                                                                           (32'h18)
`define CSRNG_REG_CMD_REQ_ACMD_LOW                                                                  (0)
`define CSRNG_REG_CMD_REQ_ACMD_MASK                                                                 (32'hf)
`define CSRNG_REG_CMD_REQ_CLEN_LOW                                                                  (4)
`define CSRNG_REG_CMD_REQ_CLEN_MASK                                                                 (32'hf0)
`define CSRNG_REG_CMD_REQ_FLAG0_LOW                                                                 (8)
`define CSRNG_REG_CMD_REQ_FLAG0_MASK                                                                (32'hf00)
`define CSRNG_REG_CMD_REQ_GLEN_LOW                                                                  (12)
`define CSRNG_REG_CMD_REQ_GLEN_MASK                                                                 (32'h1fff000)
`define CLP_CSRNG_REG_SW_CMD_STS                                                                    (32'h2000201c)
`define CSRNG_REG_SW_CMD_STS                                                                        (32'h1c)
`define CSRNG_REG_SW_CMD_STS_CMD_RDY_LOW                                                            (0)
`define CSRNG_REG_SW_CMD_STS_CMD_RDY_MASK                                                           (32'h1)
`define CSRNG_REG_SW_CMD_STS_CMD_STS_LOW                                                            (1)
`define CSRNG_REG_SW_CMD_STS_CMD_STS_MASK                                                           (32'h2)
`define CLP_CSRNG_REG_GENBITS_VLD                                                                   (32'h20002020)
`define CSRNG_REG_GENBITS_VLD                                                                       (32'h20)
`define CSRNG_REG_GENBITS_VLD_GENBITS_VLD_LOW                                                       (0)
`define CSRNG_REG_GENBITS_VLD_GENBITS_VLD_MASK                                                      (32'h1)
`define CSRNG_REG_GENBITS_VLD_GENBITS_FIPS_LOW                                                      (1)
`define CSRNG_REG_GENBITS_VLD_GENBITS_FIPS_MASK                                                     (32'h2)
`define CLP_CSRNG_REG_GENBITS                                                                       (32'h20002024)
`define CSRNG_REG_GENBITS                                                                           (32'h24)
`define CLP_CSRNG_REG_INT_STATE_NUM                                                                 (32'h20002028)
`define CSRNG_REG_INT_STATE_NUM                                                                     (32'h28)
`define CSRNG_REG_INT_STATE_NUM_INT_STATE_NUM_LOW                                                   (0)
`define CSRNG_REG_INT_STATE_NUM_INT_STATE_NUM_MASK                                                  (32'hf)
`define CLP_CSRNG_REG_INT_STATE_VAL                                                                 (32'h2000202c)
`define CSRNG_REG_INT_STATE_VAL                                                                     (32'h2c)
`define CLP_CSRNG_REG_HW_EXC_STS                                                                    (32'h20002030)
`define CSRNG_REG_HW_EXC_STS                                                                        (32'h30)
`define CSRNG_REG_HW_EXC_STS_HW_EXC_STS_LOW                                                         (0)
`define CSRNG_REG_HW_EXC_STS_HW_EXC_STS_MASK                                                        (32'hffff)
`define CLP_CSRNG_REG_RECOV_ALERT_STS                                                               (32'h20002034)
`define CSRNG_REG_RECOV_ALERT_STS                                                                   (32'h34)
`define CSRNG_REG_RECOV_ALERT_STS_ENABLE_FIELD_ALERT_LOW                                            (0)
`define CSRNG_REG_RECOV_ALERT_STS_ENABLE_FIELD_ALERT_MASK                                           (32'h1)
`define CSRNG_REG_RECOV_ALERT_STS_SW_APP_ENABLE_FIELD_ALERT_LOW                                     (1)
`define CSRNG_REG_RECOV_ALERT_STS_SW_APP_ENABLE_FIELD_ALERT_MASK                                    (32'h2)
`define CSRNG_REG_RECOV_ALERT_STS_READ_INT_STATE_FIELD_ALERT_LOW                                    (2)
`define CSRNG_REG_RECOV_ALERT_STS_READ_INT_STATE_FIELD_ALERT_MASK                                   (32'h4)
`define CSRNG_REG_RECOV_ALERT_STS_ACMD_FLAG0_FIELD_ALERT_LOW                                        (3)
`define CSRNG_REG_RECOV_ALERT_STS_ACMD_FLAG0_FIELD_ALERT_MASK                                       (32'h8)
`define CSRNG_REG_RECOV_ALERT_STS_CS_BUS_CMP_ALERT_LOW                                              (12)
`define CSRNG_REG_RECOV_ALERT_STS_CS_BUS_CMP_ALERT_MASK                                             (32'h1000)
`define CSRNG_REG_RECOV_ALERT_STS_CS_MAIN_SM_ALERT_LOW                                              (13)
`define CSRNG_REG_RECOV_ALERT_STS_CS_MAIN_SM_ALERT_MASK                                             (32'h2000)
`define CLP_CSRNG_REG_ERR_CODE                                                                      (32'h20002038)
`define CSRNG_REG_ERR_CODE                                                                          (32'h38)
`define CSRNG_REG_ERR_CODE_SFIFO_CMD_ERR_LOW                                                        (0)
`define CSRNG_REG_ERR_CODE_SFIFO_CMD_ERR_MASK                                                       (32'h1)
`define CSRNG_REG_ERR_CODE_SFIFO_GENBITS_ERR_LOW                                                    (1)
`define CSRNG_REG_ERR_CODE_SFIFO_GENBITS_ERR_MASK                                                   (32'h2)
`define CSRNG_REG_ERR_CODE_SFIFO_CMDREQ_ERR_LOW                                                     (2)
`define CSRNG_REG_ERR_CODE_SFIFO_CMDREQ_ERR_MASK                                                    (32'h4)
`define CSRNG_REG_ERR_CODE_SFIFO_RCSTAGE_ERR_LOW                                                    (3)
`define CSRNG_REG_ERR_CODE_SFIFO_RCSTAGE_ERR_MASK                                                   (32'h8)
`define CSRNG_REG_ERR_CODE_SFIFO_KEYVRC_ERR_LOW                                                     (4)
`define CSRNG_REG_ERR_CODE_SFIFO_KEYVRC_ERR_MASK                                                    (32'h10)
`define CSRNG_REG_ERR_CODE_SFIFO_UPDREQ_ERR_LOW                                                     (5)
`define CSRNG_REG_ERR_CODE_SFIFO_UPDREQ_ERR_MASK                                                    (32'h20)
`define CSRNG_REG_ERR_CODE_SFIFO_BENCREQ_ERR_LOW                                                    (6)
`define CSRNG_REG_ERR_CODE_SFIFO_BENCREQ_ERR_MASK                                                   (32'h40)
`define CSRNG_REG_ERR_CODE_SFIFO_BENCACK_ERR_LOW                                                    (7)
`define CSRNG_REG_ERR_CODE_SFIFO_BENCACK_ERR_MASK                                                   (32'h80)
`define CSRNG_REG_ERR_CODE_SFIFO_PDATA_ERR_LOW                                                      (8)
`define CSRNG_REG_ERR_CODE_SFIFO_PDATA_ERR_MASK                                                     (32'h100)
`define CSRNG_REG_ERR_CODE_SFIFO_FINAL_ERR_LOW                                                      (9)
`define CSRNG_REG_ERR_CODE_SFIFO_FINAL_ERR_MASK                                                     (32'h200)
`define CSRNG_REG_ERR_CODE_SFIFO_GBENCACK_ERR_LOW                                                   (10)
`define CSRNG_REG_ERR_CODE_SFIFO_GBENCACK_ERR_MASK                                                  (32'h400)
`define CSRNG_REG_ERR_CODE_SFIFO_GRCSTAGE_ERR_LOW                                                   (11)
`define CSRNG_REG_ERR_CODE_SFIFO_GRCSTAGE_ERR_MASK                                                  (32'h800)
`define CSRNG_REG_ERR_CODE_SFIFO_GGENREQ_ERR_LOW                                                    (12)
`define CSRNG_REG_ERR_CODE_SFIFO_GGENREQ_ERR_MASK                                                   (32'h1000)
`define CSRNG_REG_ERR_CODE_SFIFO_GADSTAGE_ERR_LOW                                                   (13)
`define CSRNG_REG_ERR_CODE_SFIFO_GADSTAGE_ERR_MASK                                                  (32'h2000)
`define CSRNG_REG_ERR_CODE_SFIFO_GGENBITS_ERR_LOW                                                   (14)
`define CSRNG_REG_ERR_CODE_SFIFO_GGENBITS_ERR_MASK                                                  (32'h4000)
`define CSRNG_REG_ERR_CODE_SFIFO_BLKENC_ERR_LOW                                                     (15)
`define CSRNG_REG_ERR_CODE_SFIFO_BLKENC_ERR_MASK                                                    (32'h8000)
`define CSRNG_REG_ERR_CODE_CMD_STAGE_SM_ERR_LOW                                                     (20)
`define CSRNG_REG_ERR_CODE_CMD_STAGE_SM_ERR_MASK                                                    (32'h100000)
`define CSRNG_REG_ERR_CODE_MAIN_SM_ERR_LOW                                                          (21)
`define CSRNG_REG_ERR_CODE_MAIN_SM_ERR_MASK                                                         (32'h200000)
`define CSRNG_REG_ERR_CODE_DRBG_GEN_SM_ERR_LOW                                                      (22)
`define CSRNG_REG_ERR_CODE_DRBG_GEN_SM_ERR_MASK                                                     (32'h400000)
`define CSRNG_REG_ERR_CODE_DRBG_UPDBE_SM_ERR_LOW                                                    (23)
`define CSRNG_REG_ERR_CODE_DRBG_UPDBE_SM_ERR_MASK                                                   (32'h800000)
`define CSRNG_REG_ERR_CODE_DRBG_UPDOB_SM_ERR_LOW                                                    (24)
`define CSRNG_REG_ERR_CODE_DRBG_UPDOB_SM_ERR_MASK                                                   (32'h1000000)
`define CSRNG_REG_ERR_CODE_AES_CIPHER_SM_ERR_LOW                                                    (25)
`define CSRNG_REG_ERR_CODE_AES_CIPHER_SM_ERR_MASK                                                   (32'h2000000)
`define CSRNG_REG_ERR_CODE_CMD_GEN_CNT_ERR_LOW                                                      (26)
`define CSRNG_REG_ERR_CODE_CMD_GEN_CNT_ERR_MASK                                                     (32'h4000000)
`define CSRNG_REG_ERR_CODE_FIFO_WRITE_ERR_LOW                                                       (28)
`define CSRNG_REG_ERR_CODE_FIFO_WRITE_ERR_MASK                                                      (32'h10000000)
`define CSRNG_REG_ERR_CODE_FIFO_READ_ERR_LOW                                                        (29)
`define CSRNG_REG_ERR_CODE_FIFO_READ_ERR_MASK                                                       (32'h20000000)
`define CSRNG_REG_ERR_CODE_FIFO_STATE_ERR_LOW                                                       (30)
`define CSRNG_REG_ERR_CODE_FIFO_STATE_ERR_MASK                                                      (32'h40000000)
`define CLP_CSRNG_REG_ERR_CODE_TEST                                                                 (32'h2000203c)
`define CSRNG_REG_ERR_CODE_TEST                                                                     (32'h3c)
`define CSRNG_REG_ERR_CODE_TEST_ERR_CODE_TEST_LOW                                                   (0)
`define CSRNG_REG_ERR_CODE_TEST_ERR_CODE_TEST_MASK                                                  (32'h1f)
`define CLP_CSRNG_REG_MAIN_SM_STATE                                                                 (32'h20002040)
`define CSRNG_REG_MAIN_SM_STATE                                                                     (32'h40)
`define CSRNG_REG_MAIN_SM_STATE_MAIN_SM_STATE_LOW                                                   (0)
`define CSRNG_REG_MAIN_SM_STATE_MAIN_SM_STATE_MASK                                                  (32'hff)
`define CLP_ENTROPY_SRC_REG_BASE_ADDR                                                               (32'h20003000)
`define CLP_ENTROPY_SRC_REG_INTERRUPT_STATE                                                         (32'h20003000)
`define ENTROPY_SRC_REG_INTERRUPT_STATE                                                             (32'h0)
`define ENTROPY_SRC_REG_INTERRUPT_STATE_ES_ENTROPY_VALID_LOW                                        (0)
`define ENTROPY_SRC_REG_INTERRUPT_STATE_ES_ENTROPY_VALID_MASK                                       (32'h1)
`define ENTROPY_SRC_REG_INTERRUPT_STATE_ES_HEALTH_TEST_FAILED_LOW                                   (1)
`define ENTROPY_SRC_REG_INTERRUPT_STATE_ES_HEALTH_TEST_FAILED_MASK                                  (32'h2)
`define ENTROPY_SRC_REG_INTERRUPT_STATE_ES_OBSERVE_FIFO_READY_LOW                                   (2)
`define ENTROPY_SRC_REG_INTERRUPT_STATE_ES_OBSERVE_FIFO_READY_MASK                                  (32'h4)
`define ENTROPY_SRC_REG_INTERRUPT_STATE_ES_FATAL_ERR_LOW                                            (3)
`define ENTROPY_SRC_REG_INTERRUPT_STATE_ES_FATAL_ERR_MASK                                           (32'h8)
`define CLP_ENTROPY_SRC_REG_INTERRUPT_ENABLE                                                        (32'h20003004)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE                                                            (32'h4)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE_ES_ENTROPY_VALID_LOW                                       (0)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE_ES_ENTROPY_VALID_MASK                                      (32'h1)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE_ES_HEALTH_TEST_FAILED_LOW                                  (1)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE_ES_HEALTH_TEST_FAILED_MASK                                 (32'h2)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE_ES_OBSERVE_FIFO_READY_LOW                                  (2)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE_ES_OBSERVE_FIFO_READY_MASK                                 (32'h4)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE_ES_FATAL_ERR_LOW                                           (3)
`define ENTROPY_SRC_REG_INTERRUPT_ENABLE_ES_FATAL_ERR_MASK                                          (32'h8)
`define CLP_ENTROPY_SRC_REG_INTERRUPT_TEST                                                          (32'h20003008)
`define ENTROPY_SRC_REG_INTERRUPT_TEST                                                              (32'h8)
`define ENTROPY_SRC_REG_INTERRUPT_TEST_ES_ENTROPY_VALID_LOW                                         (0)
`define ENTROPY_SRC_REG_INTERRUPT_TEST_ES_ENTROPY_VALID_MASK                                        (32'h1)
`define ENTROPY_SRC_REG_INTERRUPT_TEST_ES_HEALTH_TEST_FAILED_LOW                                    (1)
`define ENTROPY_SRC_REG_INTERRUPT_TEST_ES_HEALTH_TEST_FAILED_MASK                                   (32'h2)
`define ENTROPY_SRC_REG_INTERRUPT_TEST_ES_OBSERVE_FIFO_READY_LOW                                    (2)
`define ENTROPY_SRC_REG_INTERRUPT_TEST_ES_OBSERVE_FIFO_READY_MASK                                   (32'h4)
`define ENTROPY_SRC_REG_INTERRUPT_TEST_ES_FATAL_ERR_LOW                                             (3)
`define ENTROPY_SRC_REG_INTERRUPT_TEST_ES_FATAL_ERR_MASK                                            (32'h8)
`define CLP_ENTROPY_SRC_REG_ALERT_TEST                                                              (32'h2000300c)
`define ENTROPY_SRC_REG_ALERT_TEST                                                                  (32'hc)
`define ENTROPY_SRC_REG_ALERT_TEST_RECOV_ALERT_LOW                                                  (0)
`define ENTROPY_SRC_REG_ALERT_TEST_RECOV_ALERT_MASK                                                 (32'h1)
`define ENTROPY_SRC_REG_ALERT_TEST_FATAL_ALERT_LOW                                                  (1)
`define ENTROPY_SRC_REG_ALERT_TEST_FATAL_ALERT_MASK                                                 (32'h2)
`define CLP_ENTROPY_SRC_REG_ME_REGWEN                                                               (32'h20003010)
`define ENTROPY_SRC_REG_ME_REGWEN                                                                   (32'h10)
`define ENTROPY_SRC_REG_ME_REGWEN_ME_REGWEN_LOW                                                     (0)
`define ENTROPY_SRC_REG_ME_REGWEN_ME_REGWEN_MASK                                                    (32'h1)
`define CLP_ENTROPY_SRC_REG_SW_REGUPD                                                               (32'h20003014)
`define ENTROPY_SRC_REG_SW_REGUPD                                                                   (32'h14)
`define ENTROPY_SRC_REG_SW_REGUPD_SW_REGUPD_LOW                                                     (0)
`define ENTROPY_SRC_REG_SW_REGUPD_SW_REGUPD_MASK                                                    (32'h1)
`define CLP_ENTROPY_SRC_REG_REGWEN                                                                  (32'h20003018)
`define ENTROPY_SRC_REG_REGWEN                                                                      (32'h18)
`define ENTROPY_SRC_REG_REGWEN_REGWEN_LOW                                                           (0)
`define ENTROPY_SRC_REG_REGWEN_REGWEN_MASK                                                          (32'h1)
`define CLP_ENTROPY_SRC_REG_REV                                                                     (32'h2000301c)
`define ENTROPY_SRC_REG_REV                                                                         (32'h1c)
`define ENTROPY_SRC_REG_REV_ABI_REVISION_LOW                                                        (0)
`define ENTROPY_SRC_REG_REV_ABI_REVISION_MASK                                                       (32'hff)
`define ENTROPY_SRC_REG_REV_HW_REVISION_LOW                                                         (8)
`define ENTROPY_SRC_REG_REV_HW_REVISION_MASK                                                        (32'hff00)
`define ENTROPY_SRC_REG_REV_CHIP_TYPE_LOW                                                           (16)
`define ENTROPY_SRC_REG_REV_CHIP_TYPE_MASK                                                          (32'hff0000)
`define CLP_ENTROPY_SRC_REG_MODULE_ENABLE                                                           (32'h20003020)
`define ENTROPY_SRC_REG_MODULE_ENABLE                                                               (32'h20)
`define ENTROPY_SRC_REG_MODULE_ENABLE_MODULE_ENABLE_LOW                                             (0)
`define ENTROPY_SRC_REG_MODULE_ENABLE_MODULE_ENABLE_MASK                                            (32'hf)
`define CLP_ENTROPY_SRC_REG_CONF                                                                    (32'h20003024)
`define ENTROPY_SRC_REG_CONF                                                                        (32'h24)
`define ENTROPY_SRC_REG_CONF_FIPS_ENABLE_LOW                                                        (0)
`define ENTROPY_SRC_REG_CONF_FIPS_ENABLE_MASK                                                       (32'hf)
`define ENTROPY_SRC_REG_CONF_ENTROPY_DATA_REG_ENABLE_LOW                                            (4)
`define ENTROPY_SRC_REG_CONF_ENTROPY_DATA_REG_ENABLE_MASK                                           (32'hf0)
`define ENTROPY_SRC_REG_CONF_THRESHOLD_SCOPE_LOW                                                    (12)
`define ENTROPY_SRC_REG_CONF_THRESHOLD_SCOPE_MASK                                                   (32'hf000)
`define ENTROPY_SRC_REG_CONF_RNG_BIT_ENABLE_LOW                                                     (20)
`define ENTROPY_SRC_REG_CONF_RNG_BIT_ENABLE_MASK                                                    (32'hf00000)
`define ENTROPY_SRC_REG_CONF_RNG_BIT_SEL_LOW                                                        (24)
`define ENTROPY_SRC_REG_CONF_RNG_BIT_SEL_MASK                                                       (32'h3000000)
`define CLP_ENTROPY_SRC_REG_ENTROPY_CONTROL                                                         (32'h20003028)
`define ENTROPY_SRC_REG_ENTROPY_CONTROL                                                             (32'h28)
`define ENTROPY_SRC_REG_ENTROPY_CONTROL_ES_ROUTE_LOW                                                (0)
`define ENTROPY_SRC_REG_ENTROPY_CONTROL_ES_ROUTE_MASK                                               (32'hf)
`define ENTROPY_SRC_REG_ENTROPY_CONTROL_ES_TYPE_LOW                                                 (4)
`define ENTROPY_SRC_REG_ENTROPY_CONTROL_ES_TYPE_MASK                                                (32'hf0)
`define CLP_ENTROPY_SRC_REG_ENTROPY_DATA                                                            (32'h2000302c)
`define ENTROPY_SRC_REG_ENTROPY_DATA                                                                (32'h2c)
`define CLP_ENTROPY_SRC_REG_HEALTH_TEST_WINDOWS                                                     (32'h20003030)
`define ENTROPY_SRC_REG_HEALTH_TEST_WINDOWS                                                         (32'h30)
`define ENTROPY_SRC_REG_HEALTH_TEST_WINDOWS_FIPS_WINDOW_LOW                                         (0)
`define ENTROPY_SRC_REG_HEALTH_TEST_WINDOWS_FIPS_WINDOW_MASK                                        (32'hffff)
`define ENTROPY_SRC_REG_HEALTH_TEST_WINDOWS_BYPASS_WINDOW_LOW                                       (16)
`define ENTROPY_SRC_REG_HEALTH_TEST_WINDOWS_BYPASS_WINDOW_MASK                                      (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_REPCNT_THRESHOLDS                                                       (32'h20003034)
`define ENTROPY_SRC_REG_REPCNT_THRESHOLDS                                                           (32'h34)
`define ENTROPY_SRC_REG_REPCNT_THRESHOLDS_FIPS_THRESH_LOW                                           (0)
`define ENTROPY_SRC_REG_REPCNT_THRESHOLDS_FIPS_THRESH_MASK                                          (32'hffff)
`define ENTROPY_SRC_REG_REPCNT_THRESHOLDS_BYPASS_THRESH_LOW                                         (16)
`define ENTROPY_SRC_REG_REPCNT_THRESHOLDS_BYPASS_THRESH_MASK                                        (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_REPCNTS_THRESHOLDS                                                      (32'h20003038)
`define ENTROPY_SRC_REG_REPCNTS_THRESHOLDS                                                          (32'h38)
`define ENTROPY_SRC_REG_REPCNTS_THRESHOLDS_FIPS_THRESH_LOW                                          (0)
`define ENTROPY_SRC_REG_REPCNTS_THRESHOLDS_FIPS_THRESH_MASK                                         (32'hffff)
`define ENTROPY_SRC_REG_REPCNTS_THRESHOLDS_BYPASS_THRESH_LOW                                        (16)
`define ENTROPY_SRC_REG_REPCNTS_THRESHOLDS_BYPASS_THRESH_MASK                                       (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_ADAPTP_HI_THRESHOLDS                                                    (32'h2000303c)
`define ENTROPY_SRC_REG_ADAPTP_HI_THRESHOLDS                                                        (32'h3c)
`define ENTROPY_SRC_REG_ADAPTP_HI_THRESHOLDS_FIPS_THRESH_LOW                                        (0)
`define ENTROPY_SRC_REG_ADAPTP_HI_THRESHOLDS_FIPS_THRESH_MASK                                       (32'hffff)
`define ENTROPY_SRC_REG_ADAPTP_HI_THRESHOLDS_BYPASS_THRESH_LOW                                      (16)
`define ENTROPY_SRC_REG_ADAPTP_HI_THRESHOLDS_BYPASS_THRESH_MASK                                     (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_ADAPTP_LO_THRESHOLDS                                                    (32'h20003040)
`define ENTROPY_SRC_REG_ADAPTP_LO_THRESHOLDS                                                        (32'h40)
`define ENTROPY_SRC_REG_ADAPTP_LO_THRESHOLDS_FIPS_THRESH_LOW                                        (0)
`define ENTROPY_SRC_REG_ADAPTP_LO_THRESHOLDS_FIPS_THRESH_MASK                                       (32'hffff)
`define ENTROPY_SRC_REG_ADAPTP_LO_THRESHOLDS_BYPASS_THRESH_LOW                                      (16)
`define ENTROPY_SRC_REG_ADAPTP_LO_THRESHOLDS_BYPASS_THRESH_MASK                                     (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_BUCKET_THRESHOLDS                                                       (32'h20003044)
`define ENTROPY_SRC_REG_BUCKET_THRESHOLDS                                                           (32'h44)
`define ENTROPY_SRC_REG_BUCKET_THRESHOLDS_FIPS_THRESH_LOW                                           (0)
`define ENTROPY_SRC_REG_BUCKET_THRESHOLDS_FIPS_THRESH_MASK                                          (32'hffff)
`define ENTROPY_SRC_REG_BUCKET_THRESHOLDS_BYPASS_THRESH_LOW                                         (16)
`define ENTROPY_SRC_REG_BUCKET_THRESHOLDS_BYPASS_THRESH_MASK                                        (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_MARKOV_HI_THRESHOLDS                                                    (32'h20003048)
`define ENTROPY_SRC_REG_MARKOV_HI_THRESHOLDS                                                        (32'h48)
`define ENTROPY_SRC_REG_MARKOV_HI_THRESHOLDS_FIPS_THRESH_LOW                                        (0)
`define ENTROPY_SRC_REG_MARKOV_HI_THRESHOLDS_FIPS_THRESH_MASK                                       (32'hffff)
`define ENTROPY_SRC_REG_MARKOV_HI_THRESHOLDS_BYPASS_THRESH_LOW                                      (16)
`define ENTROPY_SRC_REG_MARKOV_HI_THRESHOLDS_BYPASS_THRESH_MASK                                     (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_MARKOV_LO_THRESHOLDS                                                    (32'h2000304c)
`define ENTROPY_SRC_REG_MARKOV_LO_THRESHOLDS                                                        (32'h4c)
`define ENTROPY_SRC_REG_MARKOV_LO_THRESHOLDS_FIPS_THRESH_LOW                                        (0)
`define ENTROPY_SRC_REG_MARKOV_LO_THRESHOLDS_FIPS_THRESH_MASK                                       (32'hffff)
`define ENTROPY_SRC_REG_MARKOV_LO_THRESHOLDS_BYPASS_THRESH_LOW                                      (16)
`define ENTROPY_SRC_REG_MARKOV_LO_THRESHOLDS_BYPASS_THRESH_MASK                                     (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_EXTHT_HI_THRESHOLDS                                                     (32'h20003050)
`define ENTROPY_SRC_REG_EXTHT_HI_THRESHOLDS                                                         (32'h50)
`define ENTROPY_SRC_REG_EXTHT_HI_THRESHOLDS_FIPS_THRESH_LOW                                         (0)
`define ENTROPY_SRC_REG_EXTHT_HI_THRESHOLDS_FIPS_THRESH_MASK                                        (32'hffff)
`define ENTROPY_SRC_REG_EXTHT_HI_THRESHOLDS_BYPASS_THRESH_LOW                                       (16)
`define ENTROPY_SRC_REG_EXTHT_HI_THRESHOLDS_BYPASS_THRESH_MASK                                      (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_EXTHT_LO_THRESHOLDS                                                     (32'h20003054)
`define ENTROPY_SRC_REG_EXTHT_LO_THRESHOLDS                                                         (32'h54)
`define ENTROPY_SRC_REG_EXTHT_LO_THRESHOLDS_FIPS_THRESH_LOW                                         (0)
`define ENTROPY_SRC_REG_EXTHT_LO_THRESHOLDS_FIPS_THRESH_MASK                                        (32'hffff)
`define ENTROPY_SRC_REG_EXTHT_LO_THRESHOLDS_BYPASS_THRESH_LOW                                       (16)
`define ENTROPY_SRC_REG_EXTHT_LO_THRESHOLDS_BYPASS_THRESH_MASK                                      (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_REPCNT_HI_WATERMARKS                                                    (32'h20003058)
`define ENTROPY_SRC_REG_REPCNT_HI_WATERMARKS                                                        (32'h58)
`define ENTROPY_SRC_REG_REPCNT_HI_WATERMARKS_FIPS_WATERMARK_LOW                                     (0)
`define ENTROPY_SRC_REG_REPCNT_HI_WATERMARKS_FIPS_WATERMARK_MASK                                    (32'hffff)
`define ENTROPY_SRC_REG_REPCNT_HI_WATERMARKS_BYPASS_WATERMARK_LOW                                   (16)
`define ENTROPY_SRC_REG_REPCNT_HI_WATERMARKS_BYPASS_WATERMARK_MASK                                  (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_REPCNTS_HI_WATERMARKS                                                   (32'h2000305c)
`define ENTROPY_SRC_REG_REPCNTS_HI_WATERMARKS                                                       (32'h5c)
`define ENTROPY_SRC_REG_REPCNTS_HI_WATERMARKS_FIPS_WATERMARK_LOW                                    (0)
`define ENTROPY_SRC_REG_REPCNTS_HI_WATERMARKS_FIPS_WATERMARK_MASK                                   (32'hffff)
`define ENTROPY_SRC_REG_REPCNTS_HI_WATERMARKS_BYPASS_WATERMARK_LOW                                  (16)
`define ENTROPY_SRC_REG_REPCNTS_HI_WATERMARKS_BYPASS_WATERMARK_MASK                                 (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_ADAPTP_HI_WATERMARKS                                                    (32'h20003060)
`define ENTROPY_SRC_REG_ADAPTP_HI_WATERMARKS                                                        (32'h60)
`define ENTROPY_SRC_REG_ADAPTP_HI_WATERMARKS_FIPS_WATERMARK_LOW                                     (0)
`define ENTROPY_SRC_REG_ADAPTP_HI_WATERMARKS_FIPS_WATERMARK_MASK                                    (32'hffff)
`define ENTROPY_SRC_REG_ADAPTP_HI_WATERMARKS_BYPASS_WATERMARK_LOW                                   (16)
`define ENTROPY_SRC_REG_ADAPTP_HI_WATERMARKS_BYPASS_WATERMARK_MASK                                  (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_ADAPTP_LO_WATERMARKS                                                    (32'h20003064)
`define ENTROPY_SRC_REG_ADAPTP_LO_WATERMARKS                                                        (32'h64)
`define ENTROPY_SRC_REG_ADAPTP_LO_WATERMARKS_FIPS_WATERMARK_LOW                                     (0)
`define ENTROPY_SRC_REG_ADAPTP_LO_WATERMARKS_FIPS_WATERMARK_MASK                                    (32'hffff)
`define ENTROPY_SRC_REG_ADAPTP_LO_WATERMARKS_BYPASS_WATERMARK_LOW                                   (16)
`define ENTROPY_SRC_REG_ADAPTP_LO_WATERMARKS_BYPASS_WATERMARK_MASK                                  (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_EXTHT_HI_WATERMARKS                                                     (32'h20003068)
`define ENTROPY_SRC_REG_EXTHT_HI_WATERMARKS                                                         (32'h68)
`define ENTROPY_SRC_REG_EXTHT_HI_WATERMARKS_FIPS_WATERMARK_LOW                                      (0)
`define ENTROPY_SRC_REG_EXTHT_HI_WATERMARKS_FIPS_WATERMARK_MASK                                     (32'hffff)
`define ENTROPY_SRC_REG_EXTHT_HI_WATERMARKS_BYPASS_WATERMARK_LOW                                    (16)
`define ENTROPY_SRC_REG_EXTHT_HI_WATERMARKS_BYPASS_WATERMARK_MASK                                   (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_EXTHT_LO_WATERMARKS                                                     (32'h2000306c)
`define ENTROPY_SRC_REG_EXTHT_LO_WATERMARKS                                                         (32'h6c)
`define ENTROPY_SRC_REG_EXTHT_LO_WATERMARKS_FIPS_WATERMARK_LOW                                      (0)
`define ENTROPY_SRC_REG_EXTHT_LO_WATERMARKS_FIPS_WATERMARK_MASK                                     (32'hffff)
`define ENTROPY_SRC_REG_EXTHT_LO_WATERMARKS_BYPASS_WATERMARK_LOW                                    (16)
`define ENTROPY_SRC_REG_EXTHT_LO_WATERMARKS_BYPASS_WATERMARK_MASK                                   (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_BUCKET_HI_WATERMARKS                                                    (32'h20003070)
`define ENTROPY_SRC_REG_BUCKET_HI_WATERMARKS                                                        (32'h70)
`define ENTROPY_SRC_REG_BUCKET_HI_WATERMARKS_FIPS_WATERMARK_LOW                                     (0)
`define ENTROPY_SRC_REG_BUCKET_HI_WATERMARKS_FIPS_WATERMARK_MASK                                    (32'hffff)
`define ENTROPY_SRC_REG_BUCKET_HI_WATERMARKS_BYPASS_WATERMARK_LOW                                   (16)
`define ENTROPY_SRC_REG_BUCKET_HI_WATERMARKS_BYPASS_WATERMARK_MASK                                  (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_MARKOV_HI_WATERMARKS                                                    (32'h20003074)
`define ENTROPY_SRC_REG_MARKOV_HI_WATERMARKS                                                        (32'h74)
`define ENTROPY_SRC_REG_MARKOV_HI_WATERMARKS_FIPS_WATERMARK_LOW                                     (0)
`define ENTROPY_SRC_REG_MARKOV_HI_WATERMARKS_FIPS_WATERMARK_MASK                                    (32'hffff)
`define ENTROPY_SRC_REG_MARKOV_HI_WATERMARKS_BYPASS_WATERMARK_LOW                                   (16)
`define ENTROPY_SRC_REG_MARKOV_HI_WATERMARKS_BYPASS_WATERMARK_MASK                                  (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_MARKOV_LO_WATERMARKS                                                    (32'h20003078)
`define ENTROPY_SRC_REG_MARKOV_LO_WATERMARKS                                                        (32'h78)
`define ENTROPY_SRC_REG_MARKOV_LO_WATERMARKS_FIPS_WATERMARK_LOW                                     (0)
`define ENTROPY_SRC_REG_MARKOV_LO_WATERMARKS_FIPS_WATERMARK_MASK                                    (32'hffff)
`define ENTROPY_SRC_REG_MARKOV_LO_WATERMARKS_BYPASS_WATERMARK_LOW                                   (16)
`define ENTROPY_SRC_REG_MARKOV_LO_WATERMARKS_BYPASS_WATERMARK_MASK                                  (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_REPCNT_TOTAL_FAILS                                                      (32'h2000307c)
`define ENTROPY_SRC_REG_REPCNT_TOTAL_FAILS                                                          (32'h7c)
`define CLP_ENTROPY_SRC_REG_REPCNTS_TOTAL_FAILS                                                     (32'h20003080)
`define ENTROPY_SRC_REG_REPCNTS_TOTAL_FAILS                                                         (32'h80)
`define CLP_ENTROPY_SRC_REG_ADAPTP_HI_TOTAL_FAILS                                                   (32'h20003084)
`define ENTROPY_SRC_REG_ADAPTP_HI_TOTAL_FAILS                                                       (32'h84)
`define CLP_ENTROPY_SRC_REG_ADAPTP_LO_TOTAL_FAILS                                                   (32'h20003088)
`define ENTROPY_SRC_REG_ADAPTP_LO_TOTAL_FAILS                                                       (32'h88)
`define CLP_ENTROPY_SRC_REG_BUCKET_TOTAL_FAILS                                                      (32'h2000308c)
`define ENTROPY_SRC_REG_BUCKET_TOTAL_FAILS                                                          (32'h8c)
`define CLP_ENTROPY_SRC_REG_MARKOV_HI_TOTAL_FAILS                                                   (32'h20003090)
`define ENTROPY_SRC_REG_MARKOV_HI_TOTAL_FAILS                                                       (32'h90)
`define CLP_ENTROPY_SRC_REG_MARKOV_LO_TOTAL_FAILS                                                   (32'h20003094)
`define ENTROPY_SRC_REG_MARKOV_LO_TOTAL_FAILS                                                       (32'h94)
`define CLP_ENTROPY_SRC_REG_EXTHT_HI_TOTAL_FAILS                                                    (32'h20003098)
`define ENTROPY_SRC_REG_EXTHT_HI_TOTAL_FAILS                                                        (32'h98)
`define CLP_ENTROPY_SRC_REG_EXTHT_LO_TOTAL_FAILS                                                    (32'h2000309c)
`define ENTROPY_SRC_REG_EXTHT_LO_TOTAL_FAILS                                                        (32'h9c)
`define CLP_ENTROPY_SRC_REG_ALERT_THRESHOLD                                                         (32'h200030a0)
`define ENTROPY_SRC_REG_ALERT_THRESHOLD                                                             (32'ha0)
`define ENTROPY_SRC_REG_ALERT_THRESHOLD_ALERT_THRESHOLD_LOW                                         (0)
`define ENTROPY_SRC_REG_ALERT_THRESHOLD_ALERT_THRESHOLD_MASK                                        (32'hffff)
`define ENTROPY_SRC_REG_ALERT_THRESHOLD_ALERT_THRESHOLD_INV_LOW                                     (16)
`define ENTROPY_SRC_REG_ALERT_THRESHOLD_ALERT_THRESHOLD_INV_MASK                                    (32'hffff0000)
`define CLP_ENTROPY_SRC_REG_ALERT_SUMMARY_FAIL_COUNTS                                               (32'h200030a4)
`define ENTROPY_SRC_REG_ALERT_SUMMARY_FAIL_COUNTS                                                   (32'ha4)
`define ENTROPY_SRC_REG_ALERT_SUMMARY_FAIL_COUNTS_ANY_FAIL_COUNT_LOW                                (0)
`define ENTROPY_SRC_REG_ALERT_SUMMARY_FAIL_COUNTS_ANY_FAIL_COUNT_MASK                               (32'hffff)
`define CLP_ENTROPY_SRC_REG_ALERT_FAIL_COUNTS                                                       (32'h200030a8)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS                                                           (32'ha8)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_REPCNT_FAIL_COUNT_LOW                                     (4)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_REPCNT_FAIL_COUNT_MASK                                    (32'hf0)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_ADAPTP_HI_FAIL_COUNT_LOW                                  (8)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_ADAPTP_HI_FAIL_COUNT_MASK                                 (32'hf00)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_ADAPTP_LO_FAIL_COUNT_LOW                                  (12)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_ADAPTP_LO_FAIL_COUNT_MASK                                 (32'hf000)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_BUCKET_FAIL_COUNT_LOW                                     (16)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_BUCKET_FAIL_COUNT_MASK                                    (32'hf0000)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_MARKOV_HI_FAIL_COUNT_LOW                                  (20)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_MARKOV_HI_FAIL_COUNT_MASK                                 (32'hf00000)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_MARKOV_LO_FAIL_COUNT_LOW                                  (24)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_MARKOV_LO_FAIL_COUNT_MASK                                 (32'hf000000)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_REPCNTS_FAIL_COUNT_LOW                                    (28)
`define ENTROPY_SRC_REG_ALERT_FAIL_COUNTS_REPCNTS_FAIL_COUNT_MASK                                   (32'hf0000000)
`define CLP_ENTROPY_SRC_REG_EXTHT_FAIL_COUNTS                                                       (32'h200030ac)
`define ENTROPY_SRC_REG_EXTHT_FAIL_COUNTS                                                           (32'hac)
`define ENTROPY_SRC_REG_EXTHT_FAIL_COUNTS_EXTHT_HI_FAIL_COUNT_LOW                                   (0)
`define ENTROPY_SRC_REG_EXTHT_FAIL_COUNTS_EXTHT_HI_FAIL_COUNT_MASK                                  (32'hf)
`define ENTROPY_SRC_REG_EXTHT_FAIL_COUNTS_EXTHT_LO_FAIL_COUNT_LOW                                   (4)
`define ENTROPY_SRC_REG_EXTHT_FAIL_COUNTS_EXTHT_LO_FAIL_COUNT_MASK                                  (32'hf0)
`define CLP_ENTROPY_SRC_REG_FW_OV_CONTROL                                                           (32'h200030b0)
`define ENTROPY_SRC_REG_FW_OV_CONTROL                                                               (32'hb0)
`define ENTROPY_SRC_REG_FW_OV_CONTROL_FW_OV_MODE_LOW                                                (0)
`define ENTROPY_SRC_REG_FW_OV_CONTROL_FW_OV_MODE_MASK                                               (32'hf)
`define ENTROPY_SRC_REG_FW_OV_CONTROL_FW_OV_ENTROPY_INSERT_LOW                                      (4)
`define ENTROPY_SRC_REG_FW_OV_CONTROL_FW_OV_ENTROPY_INSERT_MASK                                     (32'hf0)
`define CLP_ENTROPY_SRC_REG_FW_OV_SHA3_START                                                        (32'h200030b4)
`define ENTROPY_SRC_REG_FW_OV_SHA3_START                                                            (32'hb4)
`define ENTROPY_SRC_REG_FW_OV_SHA3_START_FW_OV_INSERT_START_LOW                                     (0)
`define ENTROPY_SRC_REG_FW_OV_SHA3_START_FW_OV_INSERT_START_MASK                                    (32'hf)
`define CLP_ENTROPY_SRC_REG_FW_OV_WR_FIFO_FULL                                                      (32'h200030b8)
`define ENTROPY_SRC_REG_FW_OV_WR_FIFO_FULL                                                          (32'hb8)
`define ENTROPY_SRC_REG_FW_OV_WR_FIFO_FULL_FW_OV_WR_FIFO_FULL_LOW                                   (0)
`define ENTROPY_SRC_REG_FW_OV_WR_FIFO_FULL_FW_OV_WR_FIFO_FULL_MASK                                  (32'h1)
`define CLP_ENTROPY_SRC_REG_FW_OV_RD_FIFO_OVERFLOW                                                  (32'h200030bc)
`define ENTROPY_SRC_REG_FW_OV_RD_FIFO_OVERFLOW                                                      (32'hbc)
`define ENTROPY_SRC_REG_FW_OV_RD_FIFO_OVERFLOW_FW_OV_RD_FIFO_OVERFLOW_LOW                           (0)
`define ENTROPY_SRC_REG_FW_OV_RD_FIFO_OVERFLOW_FW_OV_RD_FIFO_OVERFLOW_MASK                          (32'h1)
`define CLP_ENTROPY_SRC_REG_FW_OV_RD_DATA                                                           (32'h200030c0)
`define ENTROPY_SRC_REG_FW_OV_RD_DATA                                                               (32'hc0)
`define CLP_ENTROPY_SRC_REG_FW_OV_WR_DATA                                                           (32'h200030c4)
`define ENTROPY_SRC_REG_FW_OV_WR_DATA                                                               (32'hc4)
`define CLP_ENTROPY_SRC_REG_OBSERVE_FIFO_THRESH                                                     (32'h200030c8)
`define ENTROPY_SRC_REG_OBSERVE_FIFO_THRESH                                                         (32'hc8)
`define ENTROPY_SRC_REG_OBSERVE_FIFO_THRESH_OBSERVE_FIFO_THRESH_LOW                                 (0)
`define ENTROPY_SRC_REG_OBSERVE_FIFO_THRESH_OBSERVE_FIFO_THRESH_MASK                                (32'h7f)
`define CLP_ENTROPY_SRC_REG_OBSERVE_FIFO_DEPTH                                                      (32'h200030cc)
`define ENTROPY_SRC_REG_OBSERVE_FIFO_DEPTH                                                          (32'hcc)
`define ENTROPY_SRC_REG_OBSERVE_FIFO_DEPTH_OBSERVE_FIFO_DEPTH_LOW                                   (0)
`define ENTROPY_SRC_REG_OBSERVE_FIFO_DEPTH_OBSERVE_FIFO_DEPTH_MASK                                  (32'h7f)
`define CLP_ENTROPY_SRC_REG_DEBUG_STATUS                                                            (32'h200030d0)
`define ENTROPY_SRC_REG_DEBUG_STATUS                                                                (32'hd0)
`define ENTROPY_SRC_REG_DEBUG_STATUS_ENTROPY_FIFO_DEPTH_LOW                                         (0)
`define ENTROPY_SRC_REG_DEBUG_STATUS_ENTROPY_FIFO_DEPTH_MASK                                        (32'h7)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_FSM_LOW                                                   (3)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_FSM_MASK                                                  (32'h38)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_BLOCK_PR_LOW                                              (6)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_BLOCK_PR_MASK                                             (32'h40)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_SQUEEZING_LOW                                             (7)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_SQUEEZING_MASK                                            (32'h80)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_ABSORBED_LOW                                              (8)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_ABSORBED_MASK                                             (32'h100)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_ERR_LOW                                                   (9)
`define ENTROPY_SRC_REG_DEBUG_STATUS_SHA3_ERR_MASK                                                  (32'h200)
`define ENTROPY_SRC_REG_DEBUG_STATUS_MAIN_SM_IDLE_LOW                                               (16)
`define ENTROPY_SRC_REG_DEBUG_STATUS_MAIN_SM_IDLE_MASK                                              (32'h10000)
`define ENTROPY_SRC_REG_DEBUG_STATUS_MAIN_SM_BOOT_DONE_LOW                                          (17)
`define ENTROPY_SRC_REG_DEBUG_STATUS_MAIN_SM_BOOT_DONE_MASK                                         (32'h20000)
`define CLP_ENTROPY_SRC_REG_RECOV_ALERT_STS                                                         (32'h200030d4)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS                                                             (32'hd4)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_FIPS_ENABLE_FIELD_ALERT_LOW                                 (0)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_FIPS_ENABLE_FIELD_ALERT_MASK                                (32'h1)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ENTROPY_DATA_REG_EN_FIELD_ALERT_LOW                         (1)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ENTROPY_DATA_REG_EN_FIELD_ALERT_MASK                        (32'h2)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_MODULE_ENABLE_FIELD_ALERT_LOW                               (2)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_MODULE_ENABLE_FIELD_ALERT_MASK                              (32'h4)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_THRESHOLD_SCOPE_FIELD_ALERT_LOW                             (3)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_THRESHOLD_SCOPE_FIELD_ALERT_MASK                            (32'h8)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_RNG_BIT_ENABLE_FIELD_ALERT_LOW                              (5)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_RNG_BIT_ENABLE_FIELD_ALERT_MASK                             (32'h20)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_FW_OV_SHA3_START_FIELD_ALERT_LOW                            (7)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_FW_OV_SHA3_START_FIELD_ALERT_MASK                           (32'h80)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_FW_OV_MODE_FIELD_ALERT_LOW                                  (8)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_FW_OV_MODE_FIELD_ALERT_MASK                                 (32'h100)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_FW_OV_ENTROPY_INSERT_FIELD_ALERT_LOW                        (9)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_FW_OV_ENTROPY_INSERT_FIELD_ALERT_MASK                       (32'h200)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_ROUTE_FIELD_ALERT_LOW                                    (10)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_ROUTE_FIELD_ALERT_MASK                                   (32'h400)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_TYPE_FIELD_ALERT_LOW                                     (11)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_TYPE_FIELD_ALERT_MASK                                    (32'h800)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_MAIN_SM_ALERT_LOW                                        (12)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_MAIN_SM_ALERT_MASK                                       (32'h1000)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_BUS_CMP_ALERT_LOW                                        (13)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_BUS_CMP_ALERT_MASK                                       (32'h2000)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_THRESH_CFG_ALERT_LOW                                     (14)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_THRESH_CFG_ALERT_MASK                                    (32'h4000)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_FW_OV_WR_ALERT_LOW                                       (15)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_FW_OV_WR_ALERT_MASK                                      (32'h8000)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_FW_OV_DISABLE_ALERT_LOW                                  (16)
`define ENTROPY_SRC_REG_RECOV_ALERT_STS_ES_FW_OV_DISABLE_ALERT_MASK                                 (32'h10000)
`define CLP_ENTROPY_SRC_REG_ERR_CODE                                                                (32'h200030d8)
`define ENTROPY_SRC_REG_ERR_CODE                                                                    (32'hd8)
`define ENTROPY_SRC_REG_ERR_CODE_SFIFO_ESRNG_ERR_LOW                                                (0)
`define ENTROPY_SRC_REG_ERR_CODE_SFIFO_ESRNG_ERR_MASK                                               (32'h1)
`define ENTROPY_SRC_REG_ERR_CODE_SFIFO_OBSERVE_ERR_LOW                                              (1)
`define ENTROPY_SRC_REG_ERR_CODE_SFIFO_OBSERVE_ERR_MASK                                             (32'h2)
`define ENTROPY_SRC_REG_ERR_CODE_SFIFO_ESFINAL_ERR_LOW                                              (2)
`define ENTROPY_SRC_REG_ERR_CODE_SFIFO_ESFINAL_ERR_MASK                                             (32'h4)
`define ENTROPY_SRC_REG_ERR_CODE_ES_ACK_SM_ERR_LOW                                                  (20)
`define ENTROPY_SRC_REG_ERR_CODE_ES_ACK_SM_ERR_MASK                                                 (32'h100000)
`define ENTROPY_SRC_REG_ERR_CODE_ES_MAIN_SM_ERR_LOW                                                 (21)
`define ENTROPY_SRC_REG_ERR_CODE_ES_MAIN_SM_ERR_MASK                                                (32'h200000)
`define ENTROPY_SRC_REG_ERR_CODE_ES_CNTR_ERR_LOW                                                    (22)
`define ENTROPY_SRC_REG_ERR_CODE_ES_CNTR_ERR_MASK                                                   (32'h400000)
`define ENTROPY_SRC_REG_ERR_CODE_SHA3_STATE_ERR_LOW                                                 (23)
`define ENTROPY_SRC_REG_ERR_CODE_SHA3_STATE_ERR_MASK                                                (32'h800000)
`define ENTROPY_SRC_REG_ERR_CODE_SHA3_RST_STORAGE_ERR_LOW                                           (24)
`define ENTROPY_SRC_REG_ERR_CODE_SHA3_RST_STORAGE_ERR_MASK                                          (32'h1000000)
`define ENTROPY_SRC_REG_ERR_CODE_FIFO_WRITE_ERR_LOW                                                 (28)
`define ENTROPY_SRC_REG_ERR_CODE_FIFO_WRITE_ERR_MASK                                                (32'h10000000)
`define ENTROPY_SRC_REG_ERR_CODE_FIFO_READ_ERR_LOW                                                  (29)
`define ENTROPY_SRC_REG_ERR_CODE_FIFO_READ_ERR_MASK                                                 (32'h20000000)
`define ENTROPY_SRC_REG_ERR_CODE_FIFO_STATE_ERR_LOW                                                 (30)
`define ENTROPY_SRC_REG_ERR_CODE_FIFO_STATE_ERR_MASK                                                (32'h40000000)
`define CLP_ENTROPY_SRC_REG_ERR_CODE_TEST                                                           (32'h200030dc)
`define ENTROPY_SRC_REG_ERR_CODE_TEST                                                               (32'hdc)
`define ENTROPY_SRC_REG_ERR_CODE_TEST_ERR_CODE_TEST_LOW                                             (0)
`define ENTROPY_SRC_REG_ERR_CODE_TEST_ERR_CODE_TEST_MASK                                            (32'h1f)
`define CLP_ENTROPY_SRC_REG_MAIN_SM_STATE                                                           (32'h200030e0)
`define ENTROPY_SRC_REG_MAIN_SM_STATE                                                               (32'he0)
`define ENTROPY_SRC_REG_MAIN_SM_STATE_MAIN_SM_STATE_LOW                                             (0)
`define ENTROPY_SRC_REG_MAIN_SM_STATE_MAIN_SM_STATE_MASK                                            (32'h1ff)
`define CLP_MBOX_SRAM_BASE_ADDR                                                                     (32'h30000000)
`define CLP_MBOX_SRAM_END_ADDR                                                                      (32'h3001ffff)
`define CLP_MBOX_CSR_BASE_ADDR                                                                      (32'h30020000)
`define CLP_MBOX_CSR_MBOX_LOCK                                                                      (32'h30020000)
`define MBOX_CSR_MBOX_LOCK                                                                          (32'h0)
`define MBOX_CSR_MBOX_LOCK_LOCK_LOW                                                                 (0)
`define MBOX_CSR_MBOX_LOCK_LOCK_MASK                                                                (32'h1)
`define CLP_MBOX_CSR_MBOX_ID                                                                        (32'h30020004)
`define MBOX_CSR_MBOX_ID                                                                            (32'h4)
`define CLP_MBOX_CSR_MBOX_CMD                                                                       (32'h30020008)
`define MBOX_CSR_MBOX_CMD                                                                           (32'h8)
`define CLP_MBOX_CSR_MBOX_DLEN                                                                      (32'h3002000c)
`define MBOX_CSR_MBOX_DLEN                                                                          (32'hc)
`define CLP_MBOX_CSR_MBOX_DATAIN                                                                    (32'h30020010)
`define MBOX_CSR_MBOX_DATAIN                                                                        (32'h10)
`define CLP_MBOX_CSR_MBOX_DATAOUT                                                                   (32'h30020014)
`define MBOX_CSR_MBOX_DATAOUT                                                                       (32'h14)
`define CLP_MBOX_CSR_MBOX_EXECUTE                                                                   (32'h30020018)
`define MBOX_CSR_MBOX_EXECUTE                                                                       (32'h18)
`define MBOX_CSR_MBOX_EXECUTE_EXECUTE_LOW                                                           (0)
`define MBOX_CSR_MBOX_EXECUTE_EXECUTE_MASK                                                          (32'h1)
`define CLP_MBOX_CSR_MBOX_STATUS                                                                    (32'h3002001c)
`define MBOX_CSR_MBOX_STATUS                                                                        (32'h1c)
`define MBOX_CSR_MBOX_STATUS_STATUS_LOW                                                             (0)
`define MBOX_CSR_MBOX_STATUS_STATUS_MASK                                                            (32'hf)
`define MBOX_CSR_MBOX_STATUS_ECC_SINGLE_ERROR_LOW                                                   (4)
`define MBOX_CSR_MBOX_STATUS_ECC_SINGLE_ERROR_MASK                                                  (32'h10)
`define MBOX_CSR_MBOX_STATUS_ECC_DOUBLE_ERROR_LOW                                                   (5)
`define MBOX_CSR_MBOX_STATUS_ECC_DOUBLE_ERROR_MASK                                                  (32'h20)
`define MBOX_CSR_MBOX_STATUS_MBOX_FSM_PS_LOW                                                        (6)
`define MBOX_CSR_MBOX_STATUS_MBOX_FSM_PS_MASK                                                       (32'h1c0)
`define MBOX_CSR_MBOX_STATUS_SOC_HAS_LOCK_LOW                                                       (9)
`define MBOX_CSR_MBOX_STATUS_SOC_HAS_LOCK_MASK                                                      (32'h200)
`define MBOX_CSR_MBOX_STATUS_MBOX_RDPTR_LOW                                                         (10)
`define MBOX_CSR_MBOX_STATUS_MBOX_RDPTR_MASK                                                        (32'h1fffc00)
`define CLP_MBOX_CSR_MBOX_UNLOCK                                                                    (32'h30020020)
`define MBOX_CSR_MBOX_UNLOCK                                                                        (32'h20)
`define MBOX_CSR_MBOX_UNLOCK_UNLOCK_LOW                                                             (0)
`define MBOX_CSR_MBOX_UNLOCK_UNLOCK_MASK                                                            (32'h1)
`define CLP_SHA512_ACC_CSR_BASE_ADDR                                                                (32'h30021000)
`define CLP_SHA512_ACC_CSR_LOCK                                                                     (32'h30021000)
`define SHA512_ACC_CSR_LOCK                                                                         (32'h0)
`define SHA512_ACC_CSR_LOCK_LOCK_LOW                                                                (0)
`define SHA512_ACC_CSR_LOCK_LOCK_MASK                                                               (32'h1)
`define CLP_SHA512_ACC_CSR_ID                                                                       (32'h30021004)
`define SHA512_ACC_CSR_ID                                                                           (32'h4)
`define CLP_SHA512_ACC_CSR_MODE                                                                     (32'h30021008)
`define SHA512_ACC_CSR_MODE                                                                         (32'h8)
`define SHA512_ACC_CSR_MODE_MODE_LOW                                                                (0)
`define SHA512_ACC_CSR_MODE_MODE_MASK                                                               (32'h3)
`define SHA512_ACC_CSR_MODE_ENDIAN_TOGGLE_LOW                                                       (2)
`define SHA512_ACC_CSR_MODE_ENDIAN_TOGGLE_MASK                                                      (32'h4)
`define CLP_SHA512_ACC_CSR_START_ADDRESS                                                            (32'h3002100c)
`define SHA512_ACC_CSR_START_ADDRESS                                                                (32'hc)
`define CLP_SHA512_ACC_CSR_DLEN                                                                     (32'h30021010)
`define SHA512_ACC_CSR_DLEN                                                                         (32'h10)
`define CLP_SHA512_ACC_CSR_DATAIN                                                                   (32'h30021014)
`define SHA512_ACC_CSR_DATAIN                                                                       (32'h14)
`define CLP_SHA512_ACC_CSR_EXECUTE                                                                  (32'h30021018)
`define SHA512_ACC_CSR_EXECUTE                                                                      (32'h18)
`define SHA512_ACC_CSR_EXECUTE_EXECUTE_LOW                                                          (0)
`define SHA512_ACC_CSR_EXECUTE_EXECUTE_MASK                                                         (32'h1)
`define CLP_SHA512_ACC_CSR_STATUS                                                                   (32'h3002101c)
`define SHA512_ACC_CSR_STATUS                                                                       (32'h1c)
`define SHA512_ACC_CSR_STATUS_VALID_LOW                                                             (0)
`define SHA512_ACC_CSR_STATUS_VALID_MASK                                                            (32'h1)
`define SHA512_ACC_CSR_STATUS_SOC_HAS_LOCK_LOW                                                      (1)
`define SHA512_ACC_CSR_STATUS_SOC_HAS_LOCK_MASK                                                     (32'h2)
`define CLP_SHA512_ACC_CSR_DIGEST_0                                                                 (32'h30021020)
`define SHA512_ACC_CSR_DIGEST_0                                                                     (32'h20)
`define CLP_SHA512_ACC_CSR_DIGEST_1                                                                 (32'h30021024)
`define SHA512_ACC_CSR_DIGEST_1                                                                     (32'h24)
`define CLP_SHA512_ACC_CSR_DIGEST_2                                                                 (32'h30021028)
`define SHA512_ACC_CSR_DIGEST_2                                                                     (32'h28)
`define CLP_SHA512_ACC_CSR_DIGEST_3                                                                 (32'h3002102c)
`define SHA512_ACC_CSR_DIGEST_3                                                                     (32'h2c)
`define CLP_SHA512_ACC_CSR_DIGEST_4                                                                 (32'h30021030)
`define SHA512_ACC_CSR_DIGEST_4                                                                     (32'h30)
`define CLP_SHA512_ACC_CSR_DIGEST_5                                                                 (32'h30021034)
`define SHA512_ACC_CSR_DIGEST_5                                                                     (32'h34)
`define CLP_SHA512_ACC_CSR_DIGEST_6                                                                 (32'h30021038)
`define SHA512_ACC_CSR_DIGEST_6                                                                     (32'h38)
`define CLP_SHA512_ACC_CSR_DIGEST_7                                                                 (32'h3002103c)
`define SHA512_ACC_CSR_DIGEST_7                                                                     (32'h3c)
`define CLP_SHA512_ACC_CSR_DIGEST_8                                                                 (32'h30021040)
`define SHA512_ACC_CSR_DIGEST_8                                                                     (32'h40)
`define CLP_SHA512_ACC_CSR_DIGEST_9                                                                 (32'h30021044)
`define SHA512_ACC_CSR_DIGEST_9                                                                     (32'h44)
`define CLP_SHA512_ACC_CSR_DIGEST_10                                                                (32'h30021048)
`define SHA512_ACC_CSR_DIGEST_10                                                                    (32'h48)
`define CLP_SHA512_ACC_CSR_DIGEST_11                                                                (32'h3002104c)
`define SHA512_ACC_CSR_DIGEST_11                                                                    (32'h4c)
`define CLP_SHA512_ACC_CSR_DIGEST_12                                                                (32'h30021050)
`define SHA512_ACC_CSR_DIGEST_12                                                                    (32'h50)
`define CLP_SHA512_ACC_CSR_DIGEST_13                                                                (32'h30021054)
`define SHA512_ACC_CSR_DIGEST_13                                                                    (32'h54)
`define CLP_SHA512_ACC_CSR_DIGEST_14                                                                (32'h30021058)
`define SHA512_ACC_CSR_DIGEST_14                                                                    (32'h58)
`define CLP_SHA512_ACC_CSR_DIGEST_15                                                                (32'h3002105c)
`define SHA512_ACC_CSR_DIGEST_15                                                                    (32'h5c)
`define CLP_SHA512_ACC_CSR_CONTROL                                                                  (32'h30021060)
`define SHA512_ACC_CSR_CONTROL                                                                      (32'h60)
`define SHA512_ACC_CSR_CONTROL_ZEROIZE_LOW                                                          (0)
`define SHA512_ACC_CSR_CONTROL_ZEROIZE_MASK                                                         (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_START                                                      (32'h30021800)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                           (32'h30021800)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h800)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                  (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                 (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                  (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                 (32'h2)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R                                            (32'h30021804)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h804)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                  (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                 (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                  (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                 (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                  (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                 (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                  (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                 (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                            (32'h30021808)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h808)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                          (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                         (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                        (32'h3002180c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h80c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                               (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                        (32'h30021810)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h810)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                               (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                      (32'h30021814)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h814)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                           (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                          (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                           (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                          (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                           (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                          (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                           (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                          (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                      (32'h30021818)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h818)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                   (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                  (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                          (32'h3002181c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h81c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                              (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                             (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                              (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                             (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                              (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                             (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                              (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                             (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                          (32'h30021820)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h820)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                      (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                     (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                        (32'h30021900)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h900)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                        (32'h30021904)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h904)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                        (32'h30021908)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h908)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                        (32'h3002190c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h90c)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                (32'h30021980)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h980)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                   (32'h30021a00)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'ha00)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                   (32'h30021a04)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'ha04)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                   (32'h30021a08)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'ha08)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                   (32'h30021a0c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'ha0c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                           (32'h30021a10)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'ha10)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                     (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                    (32'h1)
`define CLP_AXI_DMA_REG_BASE_ADDR                                                                   (32'h30022000)
`define CLP_AXI_DMA_REG_ID                                                                          (32'h30022000)
`define AXI_DMA_REG_ID                                                                              (32'h0)
`define CLP_AXI_DMA_REG_CAP                                                                         (32'h30022004)
`define AXI_DMA_REG_CAP                                                                             (32'h4)
`define AXI_DMA_REG_CAP_FIFO_MAX_DEPTH_LOW                                                          (0)
`define AXI_DMA_REG_CAP_FIFO_MAX_DEPTH_MASK                                                         (32'hfff)
`define AXI_DMA_REG_CAP_RSVD_LOW                                                                    (12)
`define AXI_DMA_REG_CAP_RSVD_MASK                                                                   (32'hfffff000)
`define CLP_AXI_DMA_REG_CTRL                                                                        (32'h30022008)
`define AXI_DMA_REG_CTRL                                                                            (32'h8)
`define AXI_DMA_REG_CTRL_GO_LOW                                                                     (0)
`define AXI_DMA_REG_CTRL_GO_MASK                                                                    (32'h1)
`define AXI_DMA_REG_CTRL_FLUSH_LOW                                                                  (1)
`define AXI_DMA_REG_CTRL_FLUSH_MASK                                                                 (32'h2)
`define AXI_DMA_REG_CTRL_RSVD0_LOW                                                                  (2)
`define AXI_DMA_REG_CTRL_RSVD0_MASK                                                                 (32'hfffc)
`define AXI_DMA_REG_CTRL_RD_ROUTE_LOW                                                               (16)
`define AXI_DMA_REG_CTRL_RD_ROUTE_MASK                                                              (32'h30000)
`define AXI_DMA_REG_CTRL_RSVD1_LOW                                                                  (18)
`define AXI_DMA_REG_CTRL_RSVD1_MASK                                                                 (32'hc0000)
`define AXI_DMA_REG_CTRL_RD_FIXED_LOW                                                               (20)
`define AXI_DMA_REG_CTRL_RD_FIXED_MASK                                                              (32'h100000)
`define AXI_DMA_REG_CTRL_RSVD2_LOW                                                                  (21)
`define AXI_DMA_REG_CTRL_RSVD2_MASK                                                                 (32'he00000)
`define AXI_DMA_REG_CTRL_WR_ROUTE_LOW                                                               (24)
`define AXI_DMA_REG_CTRL_WR_ROUTE_MASK                                                              (32'h3000000)
`define AXI_DMA_REG_CTRL_RSVD3_LOW                                                                  (26)
`define AXI_DMA_REG_CTRL_RSVD3_MASK                                                                 (32'hc000000)
`define AXI_DMA_REG_CTRL_WR_FIXED_LOW                                                               (28)
`define AXI_DMA_REG_CTRL_WR_FIXED_MASK                                                              (32'h10000000)
`define AXI_DMA_REG_CTRL_RSVD4_LOW                                                                  (29)
`define AXI_DMA_REG_CTRL_RSVD4_MASK                                                                 (32'he0000000)
`define CLP_AXI_DMA_REG_STATUS0                                                                     (32'h3002200c)
`define AXI_DMA_REG_STATUS0                                                                         (32'hc)
`define AXI_DMA_REG_STATUS0_BUSY_LOW                                                                (0)
`define AXI_DMA_REG_STATUS0_BUSY_MASK                                                               (32'h1)
`define AXI_DMA_REG_STATUS0_ERROR_LOW                                                               (1)
`define AXI_DMA_REG_STATUS0_ERROR_MASK                                                              (32'h2)
`define AXI_DMA_REG_STATUS0_RSVD0_LOW                                                               (2)
`define AXI_DMA_REG_STATUS0_RSVD0_MASK                                                              (32'hc)
`define AXI_DMA_REG_STATUS0_FIFO_DEPTH_LOW                                                          (4)
`define AXI_DMA_REG_STATUS0_FIFO_DEPTH_MASK                                                         (32'hfff0)
`define AXI_DMA_REG_STATUS0_AXI_DMA_FSM_PS_LOW                                                      (16)
`define AXI_DMA_REG_STATUS0_AXI_DMA_FSM_PS_MASK                                                     (32'h30000)
`define AXI_DMA_REG_STATUS0_RSVD1_LOW                                                               (18)
`define AXI_DMA_REG_STATUS0_RSVD1_MASK                                                              (32'hfffc0000)
`define CLP_AXI_DMA_REG_STATUS1                                                                     (32'h30022010)
`define AXI_DMA_REG_STATUS1                                                                         (32'h10)
`define CLP_AXI_DMA_REG_SRC_ADDR_L                                                                  (32'h30022014)
`define AXI_DMA_REG_SRC_ADDR_L                                                                      (32'h14)
`define CLP_AXI_DMA_REG_SRC_ADDR_H                                                                  (32'h30022018)
`define AXI_DMA_REG_SRC_ADDR_H                                                                      (32'h18)
`define CLP_AXI_DMA_REG_DST_ADDR_L                                                                  (32'h3002201c)
`define AXI_DMA_REG_DST_ADDR_L                                                                      (32'h1c)
`define CLP_AXI_DMA_REG_DST_ADDR_H                                                                  (32'h30022020)
`define AXI_DMA_REG_DST_ADDR_H                                                                      (32'h20)
`define CLP_AXI_DMA_REG_BYTE_COUNT                                                                  (32'h30022024)
`define AXI_DMA_REG_BYTE_COUNT                                                                      (32'h24)
`define CLP_AXI_DMA_REG_BLOCK_SIZE                                                                  (32'h30022028)
`define AXI_DMA_REG_BLOCK_SIZE                                                                      (32'h28)
`define AXI_DMA_REG_BLOCK_SIZE_SIZE_LOW                                                             (0)
`define AXI_DMA_REG_BLOCK_SIZE_SIZE_MASK                                                            (32'hfff)
`define AXI_DMA_REG_BLOCK_SIZE_RSVD_LOW                                                             (12)
`define AXI_DMA_REG_BLOCK_SIZE_RSVD_MASK                                                            (32'hfffff000)
`define CLP_AXI_DMA_REG_WRITE_DATA                                                                  (32'h3002202c)
`define AXI_DMA_REG_WRITE_DATA                                                                      (32'h2c)
`define CLP_AXI_DMA_REG_READ_DATA                                                                   (32'h30022030)
`define AXI_DMA_REG_READ_DATA                                                                       (32'h30)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_START                                                         (32'h30022800)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                              (32'h30022800)
`define AXI_DMA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h800)
`define AXI_DMA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                     (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                    (32'h1)
`define AXI_DMA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                     (1)
`define AXI_DMA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                    (32'h2)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                               (32'h30022804)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h804)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_CMD_DEC_EN_LOW                              (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_CMD_DEC_EN_MASK                             (32'h1)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_AXI_RD_EN_LOW                               (1)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_AXI_RD_EN_MASK                              (32'h2)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_AXI_WR_EN_LOW                               (2)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_AXI_WR_EN_MASK                              (32'h4)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_MBOX_LOCK_EN_LOW                            (3)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_MBOX_LOCK_EN_MASK                           (32'h8)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_SHA_LOCK_EN_LOW                             (4)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_SHA_LOCK_EN_MASK                            (32'h10)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_FIFO_OFLOW_EN_LOW                           (5)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_FIFO_OFLOW_EN_MASK                          (32'h20)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_FIFO_UFLOW_EN_LOW                           (6)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_FIFO_UFLOW_EN_MASK                          (32'h40)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                               (32'h30022808)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h808)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_TXN_DONE_EN_LOW                             (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_TXN_DONE_EN_MASK                            (32'h1)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_FIFO_EMPTY_EN_LOW                           (1)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_FIFO_EMPTY_EN_MASK                          (32'h2)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_FIFO_NOT_EMPTY_EN_LOW                       (2)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_FIFO_NOT_EMPTY_EN_MASK                      (32'h4)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_FIFO_FULL_EN_LOW                            (3)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_FIFO_FULL_EN_MASK                           (32'h8)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_FIFO_NOT_FULL_EN_LOW                        (4)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_FIFO_NOT_FULL_EN_MASK                       (32'h10)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                           (32'h3002280c)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h80c)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                   (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                  (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                           (32'h30022810)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h810)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                   (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                  (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                         (32'h30022814)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h814)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_CMD_DEC_STS_LOW                       (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_CMD_DEC_STS_MASK                      (32'h1)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_AXI_RD_STS_LOW                        (1)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_AXI_RD_STS_MASK                       (32'h2)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_AXI_WR_STS_LOW                        (2)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_AXI_WR_STS_MASK                       (32'h4)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_MBOX_LOCK_STS_LOW                     (3)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_MBOX_LOCK_STS_MASK                    (32'h8)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_SHA_LOCK_STS_LOW                      (4)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_SHA_LOCK_STS_MASK                     (32'h10)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_FIFO_OFLOW_STS_LOW                    (5)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_FIFO_OFLOW_STS_MASK                   (32'h20)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_FIFO_UFLOW_STS_LOW                    (6)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_FIFO_UFLOW_STS_MASK                   (32'h40)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                         (32'h30022818)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h818)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_TXN_DONE_STS_LOW                      (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_TXN_DONE_STS_MASK                     (32'h1)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_FIFO_EMPTY_STS_LOW                    (1)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_FIFO_EMPTY_STS_MASK                   (32'h2)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_FIFO_NOT_EMPTY_STS_LOW                (2)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_FIFO_NOT_EMPTY_STS_MASK               (32'h4)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_FIFO_FULL_STS_LOW                     (3)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_FIFO_FULL_STS_MASK                    (32'h8)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_FIFO_NOT_FULL_STS_LOW                 (4)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_FIFO_NOT_FULL_STS_MASK                (32'h10)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                             (32'h3002281c)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h81c)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_CMD_DEC_TRIG_LOW                          (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_CMD_DEC_TRIG_MASK                         (32'h1)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_AXI_RD_TRIG_LOW                           (1)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_AXI_RD_TRIG_MASK                          (32'h2)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_AXI_WR_TRIG_LOW                           (2)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_AXI_WR_TRIG_MASK                          (32'h4)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_MBOX_LOCK_TRIG_LOW                        (3)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_MBOX_LOCK_TRIG_MASK                       (32'h8)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_SHA_LOCK_TRIG_LOW                         (4)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_SHA_LOCK_TRIG_MASK                        (32'h10)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_FIFO_OFLOW_TRIG_LOW                       (5)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_FIFO_OFLOW_TRIG_MASK                      (32'h20)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_FIFO_UFLOW_TRIG_LOW                       (6)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_FIFO_UFLOW_TRIG_MASK                      (32'h40)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                             (32'h30022820)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h820)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_TXN_DONE_TRIG_LOW                         (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_TXN_DONE_TRIG_MASK                        (32'h1)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_FIFO_EMPTY_TRIG_LOW                       (1)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_FIFO_EMPTY_TRIG_MASK                      (32'h2)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_FIFO_NOT_EMPTY_TRIG_LOW                   (2)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_FIFO_NOT_EMPTY_TRIG_MASK                  (32'h4)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_FIFO_FULL_TRIG_LOW                        (3)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_FIFO_FULL_TRIG_MASK                       (32'h8)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_FIFO_NOT_FULL_TRIG_LOW                    (4)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_FIFO_NOT_FULL_TRIG_MASK                   (32'h10)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_CMD_DEC_INTR_COUNT_R                                    (32'h30022900)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_CMD_DEC_INTR_COUNT_R                                        (32'h900)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_RD_INTR_COUNT_R                                     (32'h30022904)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_RD_INTR_COUNT_R                                         (32'h904)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_WR_INTR_COUNT_R                                     (32'h30022908)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_WR_INTR_COUNT_R                                         (32'h908)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_MBOX_LOCK_INTR_COUNT_R                                  (32'h3002290c)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_MBOX_LOCK_INTR_COUNT_R                                      (32'h90c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_SHA_LOCK_INTR_COUNT_R                                   (32'h30022910)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_SHA_LOCK_INTR_COUNT_R                                       (32'h910)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_OFLOW_INTR_COUNT_R                                 (32'h30022914)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_OFLOW_INTR_COUNT_R                                     (32'h914)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_UFLOW_INTR_COUNT_R                                 (32'h30022918)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_UFLOW_INTR_COUNT_R                                     (32'h918)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_TXN_DONE_INTR_COUNT_R                                   (32'h30022980)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_TXN_DONE_INTR_COUNT_R                                       (32'h980)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_EMPTY_INTR_COUNT_R                                 (32'h30022984)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_EMPTY_INTR_COUNT_R                                     (32'h984)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_EMPTY_INTR_COUNT_R                             (32'h30022988)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_EMPTY_INTR_COUNT_R                                 (32'h988)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_FULL_INTR_COUNT_R                                  (32'h3002298c)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_FULL_INTR_COUNT_R                                      (32'h98c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_FULL_INTR_COUNT_R                              (32'h30022990)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_FULL_INTR_COUNT_R                                  (32'h990)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_CMD_DEC_INTR_COUNT_INCR_R                               (32'h30022a00)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_CMD_DEC_INTR_COUNT_INCR_R                                   (32'ha00)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_CMD_DEC_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_CMD_DEC_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_RD_INTR_COUNT_INCR_R                                (32'h30022a04)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_RD_INTR_COUNT_INCR_R                                    (32'ha04)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_RD_INTR_COUNT_INCR_R_PULSE_LOW                          (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_RD_INTR_COUNT_INCR_R_PULSE_MASK                         (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_WR_INTR_COUNT_INCR_R                                (32'h30022a08)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_WR_INTR_COUNT_INCR_R                                    (32'ha08)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_WR_INTR_COUNT_INCR_R_PULSE_LOW                          (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_WR_INTR_COUNT_INCR_R_PULSE_MASK                         (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_MBOX_LOCK_INTR_COUNT_INCR_R                             (32'h30022a0c)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_MBOX_LOCK_INTR_COUNT_INCR_R                                 (32'ha0c)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_MBOX_LOCK_INTR_COUNT_INCR_R_PULSE_LOW                       (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_MBOX_LOCK_INTR_COUNT_INCR_R_PULSE_MASK                      (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_SHA_LOCK_INTR_COUNT_INCR_R                              (32'h30022a10)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_SHA_LOCK_INTR_COUNT_INCR_R                                  (32'ha10)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_SHA_LOCK_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_SHA_LOCK_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_OFLOW_INTR_COUNT_INCR_R                            (32'h30022a14)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_OFLOW_INTR_COUNT_INCR_R                                (32'ha14)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_OFLOW_INTR_COUNT_INCR_R_PULSE_LOW                      (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_OFLOW_INTR_COUNT_INCR_R_PULSE_MASK                     (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_UFLOW_INTR_COUNT_INCR_R                            (32'h30022a18)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_UFLOW_INTR_COUNT_INCR_R                                (32'ha18)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_UFLOW_INTR_COUNT_INCR_R_PULSE_LOW                      (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_UFLOW_INTR_COUNT_INCR_R_PULSE_MASK                     (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_TXN_DONE_INTR_COUNT_INCR_R                              (32'h30022a1c)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_TXN_DONE_INTR_COUNT_INCR_R                                  (32'ha1c)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_TXN_DONE_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_TXN_DONE_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_EMPTY_INTR_COUNT_INCR_R                            (32'h30022a20)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_EMPTY_INTR_COUNT_INCR_R                                (32'ha20)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_EMPTY_INTR_COUNT_INCR_R_PULSE_LOW                      (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_EMPTY_INTR_COUNT_INCR_R_PULSE_MASK                     (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_EMPTY_INTR_COUNT_INCR_R                        (32'h30022a24)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_EMPTY_INTR_COUNT_INCR_R                            (32'ha24)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_EMPTY_INTR_COUNT_INCR_R_PULSE_LOW                  (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_EMPTY_INTR_COUNT_INCR_R_PULSE_MASK                 (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_FULL_INTR_COUNT_INCR_R                             (32'h30022a28)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_FULL_INTR_COUNT_INCR_R                                 (32'ha28)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_FULL_INTR_COUNT_INCR_R_PULSE_LOW                       (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_FULL_INTR_COUNT_INCR_R_PULSE_MASK                      (32'h1)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_FULL_INTR_COUNT_INCR_R                         (32'h30022a2c)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_FULL_INTR_COUNT_INCR_R                             (32'ha2c)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_FULL_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_FULL_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)
`define CLP_SOC_IFC_REG_BASE_ADDR                                                                   (32'h30030000)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_FATAL                                                        (32'h30030000)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL                                                            (32'h0)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL_ICCM_ECC_UNC_LOW                                           (0)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL_ICCM_ECC_UNC_MASK                                          (32'h1)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL_DCCM_ECC_UNC_LOW                                           (1)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL_DCCM_ECC_UNC_MASK                                          (32'h2)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL_NMI_PIN_LOW                                                (2)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL_NMI_PIN_MASK                                               (32'h4)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL_CRYPTO_ERR_LOW                                             (3)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL_CRYPTO_ERR_MASK                                            (32'h8)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL                                                    (32'h30030004)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL                                                        (32'h4)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_PROT_NO_LOCK_LOW                                  (0)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_PROT_NO_LOCK_MASK                                 (32'h1)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_PROT_OOO_LOW                                      (1)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_PROT_OOO_MASK                                     (32'h2)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_ECC_UNC_LOW                                       (2)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_ECC_UNC_MASK                                      (32'h4)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_FATAL                                                        (32'h30030008)
`define SOC_IFC_REG_CPTRA_FW_ERROR_FATAL                                                            (32'h8)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_NON_FATAL                                                    (32'h3003000c)
`define SOC_IFC_REG_CPTRA_FW_ERROR_NON_FATAL                                                        (32'hc)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_ENC                                                          (32'h30030010)
`define SOC_IFC_REG_CPTRA_HW_ERROR_ENC                                                              (32'h10)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_ENC                                                          (32'h30030014)
`define SOC_IFC_REG_CPTRA_FW_ERROR_ENC                                                              (32'h14)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                              (32'h30030018)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                                  (32'h18)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                              (32'h3003001c)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                                  (32'h1c)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                              (32'h30030020)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                                  (32'h20)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                              (32'h30030024)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                                  (32'h24)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                              (32'h30030028)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                                  (32'h28)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                              (32'h3003002c)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                                  (32'h2c)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                              (32'h30030030)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                                  (32'h30)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                              (32'h30030034)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                                  (32'h34)
`define CLP_SOC_IFC_REG_CPTRA_BOOT_STATUS                                                           (32'h30030038)
`define SOC_IFC_REG_CPTRA_BOOT_STATUS                                                               (32'h38)
`define CLP_SOC_IFC_REG_CPTRA_FLOW_STATUS                                                           (32'h3003003c)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS                                                               (32'h3c)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_STATUS_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_STATUS_MASK                                                   (32'hffffff)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_IDEVID_CSR_READY_LOW                                          (24)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_IDEVID_CSR_READY_MASK                                         (32'h1000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_BOOT_FSM_PS_LOW                                               (25)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_BOOT_FSM_PS_MASK                                              (32'he000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FW_LOW                                              (28)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FW_MASK                                             (32'h10000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_RUNTIME_LOW                                         (29)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_RUNTIME_MASK                                        (32'h20000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FUSES_LOW                                           (30)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FUSES_MASK                                          (32'h40000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_MAILBOX_FLOW_DONE_LOW                                         (31)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_MAILBOX_FLOW_DONE_MASK                                        (32'h80000000)
`define CLP_SOC_IFC_REG_CPTRA_RESET_REASON                                                          (32'h30030040)
`define SOC_IFC_REG_CPTRA_RESET_REASON                                                              (32'h40)
`define SOC_IFC_REG_CPTRA_RESET_REASON_FW_UPD_RESET_LOW                                             (0)
`define SOC_IFC_REG_CPTRA_RESET_REASON_FW_UPD_RESET_MASK                                            (32'h1)
`define SOC_IFC_REG_CPTRA_RESET_REASON_WARM_RESET_LOW                                               (1)
`define SOC_IFC_REG_CPTRA_RESET_REASON_WARM_RESET_MASK                                              (32'h2)
`define CLP_SOC_IFC_REG_CPTRA_SECURITY_STATE                                                        (32'h30030044)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE                                                            (32'h44)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEVICE_LIFECYCLE_LOW                                       (0)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEVICE_LIFECYCLE_MASK                                      (32'h3)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEBUG_LOCKED_LOW                                           (2)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEBUG_LOCKED_MASK                                          (32'h4)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_SCAN_MODE_LOW                                              (3)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_SCAN_MODE_MASK                                             (32'h8)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_RSVD_LOW                                                   (4)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_RSVD_MASK                                                  (32'hfffffff0)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_0                                                   (32'h30030048)
`define SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_0                                                       (32'h48)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_1                                                   (32'h3003004c)
`define SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_1                                                       (32'h4c)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_2                                                   (32'h30030050)
`define SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_2                                                       (32'h50)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_3                                                   (32'h30030054)
`define SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_3                                                       (32'h54)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_4                                                   (32'h30030058)
`define SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_ID_4                                                       (32'h58)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_0                                                    (32'h3003005c)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_0                                                        (32'h5c)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_0_LOCK_LOW                                               (0)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_0_LOCK_MASK                                              (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_1                                                    (32'h30030060)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_1                                                        (32'h60)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_1_LOCK_LOW                                               (0)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_1_LOCK_MASK                                              (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_2                                                    (32'h30030064)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_2                                                        (32'h64)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_2_LOCK_LOW                                               (0)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_2_LOCK_MASK                                              (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_3                                                    (32'h30030068)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_3                                                        (32'h68)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_3_LOCK_LOW                                               (0)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_3_LOCK_MASK                                              (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_4                                                    (32'h3003006c)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_4                                                        (32'h6c)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_4_LOCK_LOW                                               (0)
`define SOC_IFC_REG_CPTRA_MBOX_AXI_ID_LOCK_4_LOCK_MASK                                              (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_VALID_AXI_ID                                                     (32'h30030070)
`define SOC_IFC_REG_CPTRA_TRNG_VALID_AXI_ID                                                         (32'h70)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_AXI_ID_LOCK                                                      (32'h30030074)
`define SOC_IFC_REG_CPTRA_TRNG_AXI_ID_LOCK                                                          (32'h74)
`define SOC_IFC_REG_CPTRA_TRNG_AXI_ID_LOCK_LOCK_LOW                                                 (0)
`define SOC_IFC_REG_CPTRA_TRNG_AXI_ID_LOCK_LOCK_MASK                                                (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_0                                                           (32'h30030078)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_0                                                               (32'h78)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_1                                                           (32'h3003007c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_1                                                               (32'h7c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_2                                                           (32'h30030080)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_2                                                               (32'h80)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_3                                                           (32'h30030084)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_3                                                               (32'h84)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_4                                                           (32'h30030088)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_4                                                               (32'h88)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_5                                                           (32'h3003008c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_5                                                               (32'h8c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_6                                                           (32'h30030090)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_6                                                               (32'h90)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_7                                                           (32'h30030094)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_7                                                               (32'h94)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_8                                                           (32'h30030098)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_8                                                               (32'h98)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_9                                                           (32'h3003009c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_9                                                               (32'h9c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_10                                                          (32'h300300a0)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_10                                                              (32'ha0)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_11                                                          (32'h300300a4)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_11                                                              (32'ha4)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_CTRL                                                             (32'h300300a8)
`define SOC_IFC_REG_CPTRA_TRNG_CTRL                                                                 (32'ha8)
`define SOC_IFC_REG_CPTRA_TRNG_CTRL_CLEAR_LOW                                                       (0)
`define SOC_IFC_REG_CPTRA_TRNG_CTRL_CLEAR_MASK                                                      (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_STATUS                                                           (32'h300300ac)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS                                                               (32'hac)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_REQ_LOW                                                  (0)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_REQ_MASK                                                 (32'h1)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_WR_DONE_LOW                                              (1)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_WR_DONE_MASK                                             (32'h2)
`define CLP_SOC_IFC_REG_CPTRA_FUSE_WR_DONE                                                          (32'h300300b0)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE                                                              (32'hb0)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE_DONE_LOW                                                     (0)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE_DONE_MASK                                                    (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TIMER_CONFIG                                                          (32'h300300b4)
`define SOC_IFC_REG_CPTRA_TIMER_CONFIG                                                              (32'hb4)
`define CLP_SOC_IFC_REG_CPTRA_BOOTFSM_GO                                                            (32'h300300b8)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO                                                                (32'hb8)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO_GO_LOW                                                         (0)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO_GO_MASK                                                        (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG                                                 (32'h300300bc)
`define SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG                                                     (32'hbc)
`define CLP_SOC_IFC_REG_CPTRA_CLK_GATING_EN                                                         (32'h300300c0)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN                                                             (32'hc0)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN_CLK_GATING_EN_LOW                                           (0)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN_CLK_GATING_EN_MASK                                          (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_0                                                 (32'h300300c4)
`define SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_0                                                     (32'hc4)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_1                                                 (32'h300300c8)
`define SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_1                                                     (32'hc8)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                                (32'h300300cc)
`define SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                                    (32'hcc)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                                (32'h300300d0)
`define SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                                    (32'hd0)
`define CLP_SOC_IFC_REG_CPTRA_HW_REV_ID                                                             (32'h300300d4)
`define SOC_IFC_REG_CPTRA_HW_REV_ID                                                                 (32'hd4)
`define SOC_IFC_REG_CPTRA_HW_REV_ID_CPTRA_GENERATION_LOW                                            (0)
`define SOC_IFC_REG_CPTRA_HW_REV_ID_CPTRA_GENERATION_MASK                                           (32'hffff)
`define SOC_IFC_REG_CPTRA_HW_REV_ID_SOC_STEPPING_ID_LOW                                             (16)
`define SOC_IFC_REG_CPTRA_HW_REV_ID_SOC_STEPPING_ID_MASK                                            (32'hffff0000)
`define CLP_SOC_IFC_REG_CPTRA_FW_REV_ID_0                                                           (32'h300300d8)
`define SOC_IFC_REG_CPTRA_FW_REV_ID_0                                                               (32'hd8)
`define CLP_SOC_IFC_REG_CPTRA_FW_REV_ID_1                                                           (32'h300300dc)
`define SOC_IFC_REG_CPTRA_FW_REV_ID_1                                                               (32'hdc)
`define CLP_SOC_IFC_REG_CPTRA_HW_CONFIG                                                             (32'h300300e0)
`define SOC_IFC_REG_CPTRA_HW_CONFIG                                                                 (32'he0)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_ITRNG_EN_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_ITRNG_EN_MASK                                                   (32'h1)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_QSPI_EN_LOW                                                     (1)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_QSPI_EN_MASK                                                    (32'h2)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_I3C_EN_LOW                                                      (2)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_I3C_EN_MASK                                                     (32'h4)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_UART_EN_LOW                                                     (3)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_UART_EN_MASK                                                    (32'h8)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_LMS_ACC_EN_LOW                                                  (4)
`define SOC_IFC_REG_CPTRA_HW_CONFIG_LMS_ACC_EN_MASK                                                 (32'h10)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER1_EN                                                         (32'h300300e4)
`define SOC_IFC_REG_CPTRA_WDT_TIMER1_EN                                                             (32'he4)
`define SOC_IFC_REG_CPTRA_WDT_TIMER1_EN_TIMER1_EN_LOW                                               (0)
`define SOC_IFC_REG_CPTRA_WDT_TIMER1_EN_TIMER1_EN_MASK                                              (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER1_CTRL                                                       (32'h300300e8)
`define SOC_IFC_REG_CPTRA_WDT_TIMER1_CTRL                                                           (32'he8)
`define SOC_IFC_REG_CPTRA_WDT_TIMER1_CTRL_TIMER1_RESTART_LOW                                        (0)
`define SOC_IFC_REG_CPTRA_WDT_TIMER1_CTRL_TIMER1_RESTART_MASK                                       (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_0                                           (32'h300300ec)
`define SOC_IFC_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_0                                               (32'hec)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_1                                           (32'h300300f0)
`define SOC_IFC_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_1                                               (32'hf0)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER2_EN                                                         (32'h300300f4)
`define SOC_IFC_REG_CPTRA_WDT_TIMER2_EN                                                             (32'hf4)
`define SOC_IFC_REG_CPTRA_WDT_TIMER2_EN_TIMER2_EN_LOW                                               (0)
`define SOC_IFC_REG_CPTRA_WDT_TIMER2_EN_TIMER2_EN_MASK                                              (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER2_CTRL                                                       (32'h300300f8)
`define SOC_IFC_REG_CPTRA_WDT_TIMER2_CTRL                                                           (32'hf8)
`define SOC_IFC_REG_CPTRA_WDT_TIMER2_CTRL_TIMER2_RESTART_LOW                                        (0)
`define SOC_IFC_REG_CPTRA_WDT_TIMER2_CTRL_TIMER2_RESTART_MASK                                       (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_0                                           (32'h300300fc)
`define SOC_IFC_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_0                                               (32'hfc)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_1                                           (32'h30030100)
`define SOC_IFC_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_1                                               (32'h100)
`define CLP_SOC_IFC_REG_CPTRA_WDT_STATUS                                                            (32'h30030104)
`define SOC_IFC_REG_CPTRA_WDT_STATUS                                                                (32'h104)
`define SOC_IFC_REG_CPTRA_WDT_STATUS_T1_TIMEOUT_LOW                                                 (0)
`define SOC_IFC_REG_CPTRA_WDT_STATUS_T1_TIMEOUT_MASK                                                (32'h1)
`define SOC_IFC_REG_CPTRA_WDT_STATUS_T2_TIMEOUT_LOW                                                 (1)
`define SOC_IFC_REG_CPTRA_WDT_STATUS_T2_TIMEOUT_MASK                                                (32'h2)
`define CLP_SOC_IFC_REG_CPTRA_FUSE_VALID_AXI_ID                                                     (32'h30030108)
`define SOC_IFC_REG_CPTRA_FUSE_VALID_AXI_ID                                                         (32'h108)
`define CLP_SOC_IFC_REG_CPTRA_FUSE_AXI_ID_LOCK                                                      (32'h3003010c)
`define SOC_IFC_REG_CPTRA_FUSE_AXI_ID_LOCK                                                          (32'h10c)
`define SOC_IFC_REG_CPTRA_FUSE_AXI_ID_LOCK_LOCK_LOW                                                 (0)
`define SOC_IFC_REG_CPTRA_FUSE_AXI_ID_LOCK_LOCK_MASK                                                (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_WDT_CFG_0                                                             (32'h30030110)
`define SOC_IFC_REG_CPTRA_WDT_CFG_0                                                                 (32'h110)
`define CLP_SOC_IFC_REG_CPTRA_WDT_CFG_1                                                             (32'h30030114)
`define SOC_IFC_REG_CPTRA_WDT_CFG_1                                                                 (32'h114)
`define CLP_SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0                                                (32'h30030118)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0                                                    (32'h118)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0_LOW_THRESHOLD_LOW                                  (0)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0_LOW_THRESHOLD_MASK                                 (32'hffff)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0_HIGH_THRESHOLD_LOW                                 (16)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0_HIGH_THRESHOLD_MASK                                (32'hffff0000)
`define CLP_SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1                                                (32'h3003011c)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1                                                    (32'h11c)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1_REPETITION_COUNT_LOW                               (0)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1_REPETITION_COUNT_MASK                              (32'hffff)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1_RSVD_LOW                                           (16)
`define SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1_RSVD_MASK                                          (32'hffff0000)
`define CLP_SOC_IFC_REG_CPTRA_RSVD_REG_0                                                            (32'h30030120)
`define SOC_IFC_REG_CPTRA_RSVD_REG_0                                                                (32'h120)
`define CLP_SOC_IFC_REG_CPTRA_RSVD_REG_1                                                            (32'h30030124)
`define SOC_IFC_REG_CPTRA_RSVD_REG_1                                                                (32'h124)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_0                                                             (32'h30030200)
`define SOC_IFC_REG_FUSE_UDS_SEED_0                                                                 (32'h200)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_1                                                             (32'h30030204)
`define SOC_IFC_REG_FUSE_UDS_SEED_1                                                                 (32'h204)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_2                                                             (32'h30030208)
`define SOC_IFC_REG_FUSE_UDS_SEED_2                                                                 (32'h208)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_3                                                             (32'h3003020c)
`define SOC_IFC_REG_FUSE_UDS_SEED_3                                                                 (32'h20c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_4                                                             (32'h30030210)
`define SOC_IFC_REG_FUSE_UDS_SEED_4                                                                 (32'h210)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_5                                                             (32'h30030214)
`define SOC_IFC_REG_FUSE_UDS_SEED_5                                                                 (32'h214)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_6                                                             (32'h30030218)
`define SOC_IFC_REG_FUSE_UDS_SEED_6                                                                 (32'h218)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_7                                                             (32'h3003021c)
`define SOC_IFC_REG_FUSE_UDS_SEED_7                                                                 (32'h21c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_8                                                             (32'h30030220)
`define SOC_IFC_REG_FUSE_UDS_SEED_8                                                                 (32'h220)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_9                                                             (32'h30030224)
`define SOC_IFC_REG_FUSE_UDS_SEED_9                                                                 (32'h224)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_10                                                            (32'h30030228)
`define SOC_IFC_REG_FUSE_UDS_SEED_10                                                                (32'h228)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_11                                                            (32'h3003022c)
`define SOC_IFC_REG_FUSE_UDS_SEED_11                                                                (32'h22c)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_0                                                        (32'h30030230)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_0                                                            (32'h230)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_1                                                        (32'h30030234)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_1                                                            (32'h234)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_2                                                        (32'h30030238)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_2                                                            (32'h238)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_3                                                        (32'h3003023c)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_3                                                            (32'h23c)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_4                                                        (32'h30030240)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_4                                                            (32'h240)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_5                                                        (32'h30030244)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_5                                                            (32'h244)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_6                                                        (32'h30030248)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_6                                                            (32'h248)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_7                                                        (32'h3003024c)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_7                                                            (32'h24c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_0                                                 (32'h30030250)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_0                                                     (32'h250)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_1                                                 (32'h30030254)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_1                                                     (32'h254)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_2                                                 (32'h30030258)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_2                                                     (32'h258)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_3                                                 (32'h3003025c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_3                                                     (32'h25c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_4                                                 (32'h30030260)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_4                                                     (32'h260)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_5                                                 (32'h30030264)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_5                                                     (32'h264)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_6                                                 (32'h30030268)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_6                                                     (32'h268)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_7                                                 (32'h3003026c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_7                                                     (32'h26c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_8                                                 (32'h30030270)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_8                                                     (32'h270)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_9                                                 (32'h30030274)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_9                                                     (32'h274)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_10                                                (32'h30030278)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_10                                                    (32'h278)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_11                                                (32'h3003027c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_11                                                    (32'h27c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK                                              (32'h30030280)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK                                                  (32'h280)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK_MASK_LOW                                         (0)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK_MASK_MASK                                        (32'hf)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_0                                                        (32'h30030284)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_0                                                            (32'h284)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_1                                                        (32'h30030288)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_1                                                            (32'h288)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_2                                                        (32'h3003028c)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_2                                                            (32'h28c)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_3                                                        (32'h30030290)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_3                                                            (32'h290)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_4                                                        (32'h30030294)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_4                                                            (32'h294)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_5                                                        (32'h30030298)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_5                                                            (32'h298)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_6                                                        (32'h3003029c)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_6                                                            (32'h29c)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_7                                                        (32'h300302a0)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_7                                                            (32'h2a0)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_8                                                        (32'h300302a4)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_8                                                            (32'h2a4)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_9                                                        (32'h300302a8)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_9                                                            (32'h2a8)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_10                                                       (32'h300302ac)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_10                                                           (32'h2ac)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_11                                                       (32'h300302b0)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_11                                                           (32'h2b0)
`define CLP_SOC_IFC_REG_FUSE_FMC_KEY_MANIFEST_SVN                                                   (32'h300302b4)
`define SOC_IFC_REG_FUSE_FMC_KEY_MANIFEST_SVN                                                       (32'h2b4)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_0                                                          (32'h300302b8)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_0                                                              (32'h2b8)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_1                                                          (32'h300302bc)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_1                                                              (32'h2bc)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_2                                                          (32'h300302c0)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_2                                                              (32'h2c0)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_3                                                          (32'h300302c4)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_3                                                              (32'h2c4)
`define CLP_SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE                                                  (32'h300302c8)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE                                                      (32'h2c8)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE_DIS_LOW                                              (0)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE_DIS_MASK                                             (32'h1)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_0                                                     (32'h300302cc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_0                                                         (32'h2cc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_1                                                     (32'h300302d0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_1                                                         (32'h2d0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_2                                                     (32'h300302d4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_2                                                         (32'h2d4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_3                                                     (32'h300302d8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_3                                                         (32'h2d8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_4                                                     (32'h300302dc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_4                                                         (32'h2dc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_5                                                     (32'h300302e0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_5                                                         (32'h2e0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6                                                     (32'h300302e4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6                                                         (32'h2e4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7                                                     (32'h300302e8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7                                                         (32'h2e8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8                                                     (32'h300302ec)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8                                                         (32'h2ec)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9                                                     (32'h300302f0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9                                                         (32'h2f0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10                                                    (32'h300302f4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10                                                        (32'h2f4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_11                                                    (32'h300302f8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_11                                                        (32'h2f8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_12                                                    (32'h300302fc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_12                                                        (32'h2fc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_13                                                    (32'h30030300)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_13                                                        (32'h300)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_14                                                    (32'h30030304)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_14                                                        (32'h304)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_15                                                    (32'h30030308)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_15                                                        (32'h308)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_16                                                    (32'h3003030c)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_16                                                        (32'h30c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_17                                                    (32'h30030310)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_17                                                        (32'h310)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_18                                                    (32'h30030314)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_18                                                        (32'h314)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_19                                                    (32'h30030318)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_19                                                        (32'h318)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_20                                                    (32'h3003031c)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_20                                                        (32'h31c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_21                                                    (32'h30030320)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_21                                                        (32'h320)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_22                                                    (32'h30030324)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_22                                                        (32'h324)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_23                                                    (32'h30030328)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_23                                                        (32'h328)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                                  (32'h3003032c)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                                      (32'h32c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                                  (32'h30030330)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                                      (32'h330)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                                  (32'h30030334)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                                      (32'h334)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                                  (32'h30030338)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                                      (32'h338)
`define CLP_SOC_IFC_REG_FUSE_LIFE_CYCLE                                                             (32'h3003033c)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE                                                                 (32'h33c)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE_LIFE_CYCLE_LOW                                                  (0)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE_LIFE_CYCLE_MASK                                                 (32'h3)
`define CLP_SOC_IFC_REG_FUSE_LMS_VERIFY                                                             (32'h30030340)
`define SOC_IFC_REG_FUSE_LMS_VERIFY                                                                 (32'h340)
`define SOC_IFC_REG_FUSE_LMS_VERIFY_LMS_VERIFY_LOW                                                  (0)
`define SOC_IFC_REG_FUSE_LMS_VERIFY_LMS_VERIFY_MASK                                                 (32'h1)
`define CLP_SOC_IFC_REG_FUSE_LMS_REVOCATION                                                         (32'h30030344)
`define SOC_IFC_REG_FUSE_LMS_REVOCATION                                                             (32'h344)
`define CLP_SOC_IFC_REG_FUSE_SOC_STEPPING_ID                                                        (32'h30030348)
`define SOC_IFC_REG_FUSE_SOC_STEPPING_ID                                                            (32'h348)
`define SOC_IFC_REG_FUSE_SOC_STEPPING_ID_SOC_STEPPING_ID_LOW                                        (0)
`define SOC_IFC_REG_FUSE_SOC_STEPPING_ID_SOC_STEPPING_ID_MASK                                       (32'hffff)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_0                                                          (32'h30030600)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_0                                                              (32'h600)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_1                                                          (32'h30030604)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_1                                                              (32'h604)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_2                                                          (32'h30030608)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_2                                                              (32'h608)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_3                                                          (32'h3003060c)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_3                                                              (32'h60c)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_4                                                          (32'h30030610)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_4                                                              (32'h610)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_5                                                          (32'h30030614)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_5                                                              (32'h614)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_6                                                          (32'h30030618)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_6                                                              (32'h618)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_7                                                          (32'h3003061c)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_7                                                              (32'h61c)
`define CLP_SOC_IFC_REG_INTERNAL_ICCM_LOCK                                                          (32'h30030620)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK                                                              (32'h620)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK_LOCK_LOW                                                     (0)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK_LOCK_MASK                                                    (32'h1)
`define CLP_SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET                                                    (32'h30030624)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET                                                        (32'h624)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_CORE_RST_LOW                                           (0)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_CORE_RST_MASK                                          (32'h1)
`define CLP_SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES                                        (32'h30030628)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES                                            (32'h628)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES_WAIT_CYCLES_LOW                            (0)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES_WAIT_CYCLES_MASK                           (32'hff)
`define CLP_SOC_IFC_REG_INTERNAL_NMI_VECTOR                                                         (32'h3003062c)
`define SOC_IFC_REG_INTERNAL_NMI_VECTOR                                                             (32'h62c)
`define CLP_SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK                                                (32'h30030630)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK                                                    (32'h630)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_ICCM_ECC_UNC_LOW                              (0)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_ICCM_ECC_UNC_MASK                             (32'h1)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_DCCM_ECC_UNC_LOW                              (1)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_DCCM_ECC_UNC_MASK                             (32'h2)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_NMI_PIN_LOW                                   (2)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_NMI_PIN_MASK                                  (32'h4)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_CRYPTO_ERR_LOW                                (3)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK_MASK_CRYPTO_ERR_MASK                               (32'h8)
`define CLP_SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK                                            (32'h30030634)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK                                                (32'h634)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK_MASK_MBOX_PROT_NO_LOCK_LOW                     (0)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK_MASK_MBOX_PROT_NO_LOCK_MASK                    (32'h1)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK_MASK_MBOX_PROT_OOO_LOW                         (1)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK_MASK_MBOX_PROT_OOO_MASK                        (32'h2)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK_MASK_MBOX_ECC_UNC_LOW                          (2)
`define SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK_MASK_MBOX_ECC_UNC_MASK                         (32'h4)
`define CLP_SOC_IFC_REG_INTERNAL_FW_ERROR_FATAL_MASK                                                (32'h30030638)
`define SOC_IFC_REG_INTERNAL_FW_ERROR_FATAL_MASK                                                    (32'h638)
`define CLP_SOC_IFC_REG_INTERNAL_FW_ERROR_NON_FATAL_MASK                                            (32'h3003063c)
`define SOC_IFC_REG_INTERNAL_FW_ERROR_NON_FATAL_MASK                                                (32'h63c)
`define CLP_SOC_IFC_REG_INTERNAL_RV_MTIME_L                                                         (32'h30030640)
`define SOC_IFC_REG_INTERNAL_RV_MTIME_L                                                             (32'h640)
`define CLP_SOC_IFC_REG_INTERNAL_RV_MTIME_H                                                         (32'h30030644)
`define SOC_IFC_REG_INTERNAL_RV_MTIME_H                                                             (32'h644)
`define CLP_SOC_IFC_REG_INTERNAL_RV_MTIMECMP_L                                                      (32'h30030648)
`define SOC_IFC_REG_INTERNAL_RV_MTIMECMP_L                                                          (32'h648)
`define CLP_SOC_IFC_REG_INTERNAL_RV_MTIMECMP_H                                                      (32'h3003064c)
`define SOC_IFC_REG_INTERNAL_RV_MTIMECMP_H                                                          (32'h64c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_START                                                         (32'h30030800)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                              (32'h30030800)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h800)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                     (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                    (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                     (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                    (32'h2)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                               (32'h30030804)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h804)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_LOW                             (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_MASK                            (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INV_DEV_EN_LOW                              (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INV_DEV_EN_MASK                             (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_CMD_FAIL_EN_LOW                             (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_CMD_FAIL_EN_MASK                            (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_BAD_FUSE_EN_LOW                             (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_BAD_FUSE_EN_MASK                            (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_ICCM_BLOCKED_EN_LOW                         (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_ICCM_BLOCKED_EN_MASK                        (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_MBOX_ECC_UNC_EN_LOW                         (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_MBOX_ECC_UNC_EN_MASK                        (32'h20)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_WDT_TIMER1_TIMEOUT_EN_LOW                   (6)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_WDT_TIMER1_TIMEOUT_EN_MASK                  (32'h40)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_WDT_TIMER2_TIMEOUT_EN_LOW                   (7)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_WDT_TIMER2_TIMEOUT_EN_MASK                  (32'h80)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                               (32'h30030808)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h808)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_AVAIL_EN_LOW                            (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_AVAIL_EN_MASK                           (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_MBOX_ECC_COR_EN_LOW                         (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_MBOX_ECC_COR_EN_MASK                        (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_DEBUG_LOCKED_EN_LOW                         (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_DEBUG_LOCKED_EN_MASK                        (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_SCAN_MODE_EN_LOW                            (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_SCAN_MODE_EN_MASK                           (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_SOC_REQ_LOCK_EN_LOW                         (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_SOC_REQ_LOCK_EN_MASK                        (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_GEN_IN_TOGGLE_EN_LOW                        (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_GEN_IN_TOGGLE_EN_MASK                       (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                           (32'h3003080c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h80c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                   (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                  (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                           (32'h30030810)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h810)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                   (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                  (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                         (32'h30030814)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h814)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_LOW                      (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_MASK                     (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INV_DEV_STS_LOW                       (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INV_DEV_STS_MASK                      (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_CMD_FAIL_STS_LOW                      (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_CMD_FAIL_STS_MASK                     (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_BAD_FUSE_STS_LOW                      (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_BAD_FUSE_STS_MASK                     (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_ICCM_BLOCKED_STS_LOW                  (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_ICCM_BLOCKED_STS_MASK                 (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_MBOX_ECC_UNC_STS_LOW                  (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_MBOX_ECC_UNC_STS_MASK                 (32'h20)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_WDT_TIMER1_TIMEOUT_STS_LOW            (6)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_WDT_TIMER1_TIMEOUT_STS_MASK           (32'h40)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_WDT_TIMER2_TIMEOUT_STS_LOW            (7)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_WDT_TIMER2_TIMEOUT_STS_MASK           (32'h80)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                         (32'h30030818)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h818)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_AVAIL_STS_LOW                     (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_AVAIL_STS_MASK                    (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_MBOX_ECC_COR_STS_LOW                  (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_MBOX_ECC_COR_STS_MASK                 (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_DEBUG_LOCKED_STS_LOW                  (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_DEBUG_LOCKED_STS_MASK                 (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_SCAN_MODE_STS_LOW                     (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_SCAN_MODE_STS_MASK                    (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_SOC_REQ_LOCK_STS_LOW                  (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_SOC_REQ_LOCK_STS_MASK                 (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_GEN_IN_TOGGLE_STS_LOW                 (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_GEN_IN_TOGGLE_STS_MASK                (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                             (32'h3003081c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h81c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_LOW                         (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_MASK                        (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INV_DEV_TRIG_LOW                          (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INV_DEV_TRIG_MASK                         (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_CMD_FAIL_TRIG_LOW                         (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_CMD_FAIL_TRIG_MASK                        (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_BAD_FUSE_TRIG_LOW                         (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_BAD_FUSE_TRIG_MASK                        (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_ICCM_BLOCKED_TRIG_LOW                     (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_ICCM_BLOCKED_TRIG_MASK                    (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_MBOX_ECC_UNC_TRIG_LOW                     (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_MBOX_ECC_UNC_TRIG_MASK                    (32'h20)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_WDT_TIMER1_TIMEOUT_TRIG_LOW               (6)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_WDT_TIMER1_TIMEOUT_TRIG_MASK              (32'h40)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_WDT_TIMER2_TIMEOUT_TRIG_LOW               (7)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_WDT_TIMER2_TIMEOUT_TRIG_MASK              (32'h80)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                             (32'h30030820)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h820)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_AVAIL_TRIG_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_AVAIL_TRIG_MASK                       (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_MBOX_ECC_COR_TRIG_LOW                     (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_MBOX_ECC_COR_TRIG_MASK                    (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_DEBUG_LOCKED_TRIG_LOW                     (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_DEBUG_LOCKED_TRIG_MASK                    (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_SCAN_MODE_TRIG_LOW                        (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_SCAN_MODE_TRIG_MASK                       (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_SOC_REQ_LOCK_TRIG_LOW                     (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_SOC_REQ_LOCK_TRIG_MASK                    (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_GEN_IN_TOGGLE_TRIG_LOW                    (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_GEN_IN_TOGGLE_TRIG_MASK                   (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                   (32'h30030900)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h900)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_R                                    (32'h30030904)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_R                                        (32'h904)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_R                                   (32'h30030908)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_R                                       (32'h908)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_R                                   (32'h3003090c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_R                                       (32'h90c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_R                               (32'h30030910)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_R                                   (32'h910)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_R                               (32'h30030914)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_R                                   (32'h914)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_R                         (32'h30030918)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_R                             (32'h918)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_R                         (32'h3003091c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_R                             (32'h91c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_R                                  (32'h30030980)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_R                                      (32'h980)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_R                               (32'h30030984)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_R                                   (32'h984)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                               (32'h30030988)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                                   (32'h988)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_R                                  (32'h3003098c)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_R                                      (32'h98c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SOC_REQ_LOCK_INTR_COUNT_R                               (32'h30030990)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SOC_REQ_LOCK_INTR_COUNT_R                                   (32'h990)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_R                              (32'h30030994)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_R                                  (32'h994)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                              (32'h30030a00)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'ha00)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R                               (32'h30030a04)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R                                   (32'ha04)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R                              (32'h30030a08)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R                                  (32'ha08)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R                              (32'h30030a0c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R                                  (32'ha0c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R                          (32'h30030a10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R                              (32'ha10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R                          (32'h30030a14)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R                              (32'ha14)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R                    (32'h30030a18)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R                        (32'ha18)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R_PULSE_LOW              (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R_PULSE_MASK             (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R                    (32'h30030a1c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R                        (32'ha1c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R_PULSE_LOW              (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R_PULSE_MASK             (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R                             (32'h30030a20)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R                                 (32'ha20)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R_PULSE_LOW                       (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R_PULSE_MASK                      (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R                          (32'h30030a24)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R                              (32'ha24)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                          (32'h30030a28)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                              (32'ha28)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_INCR_R                             (32'h30030a2c)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_INCR_R                                 (32'ha2c)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_INCR_R_PULSE_LOW                       (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_INCR_R_PULSE_MASK                      (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SOC_REQ_LOCK_INTR_COUNT_INCR_R                          (32'h30030a30)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SOC_REQ_LOCK_INTR_COUNT_INCR_R                              (32'ha30)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SOC_REQ_LOCK_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SOC_REQ_LOCK_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_INCR_R                         (32'h30030a34)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_INCR_R                             (32'ha34)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_INCR_R_PULSE_LOW                   (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_INCR_R_PULSE_MASK                  (32'h1)


`endif