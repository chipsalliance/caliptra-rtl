// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package caliptra_prim_sparse_fsm_pkg;
  typedef enum logic {Idle, Done} state_t;
endpackage : caliptra_prim_sparse_fsm_pkg
