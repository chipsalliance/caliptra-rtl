// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// Generated by PeakRDL-regblock - A free and open-source SystemVerilog generator
//  https://github.com/SystemRDL/PeakRDL-regblock

module ecc_reg (
        input wire clk,
        input wire rst,

        input wire s_cpuif_req,
        input wire s_cpuif_req_is_wr,
        input wire [10:0] s_cpuif_addr,
        input wire [31:0] s_cpuif_wr_data,
        output wire s_cpuif_req_stall_wr,
        output wire s_cpuif_req_stall_rd,
        output wire s_cpuif_rd_ack,
        output wire s_cpuif_rd_err,
        output wire [31:0] s_cpuif_rd_data,
        output wire s_cpuif_wr_ack,
        output wire s_cpuif_wr_err,

        input ecc_reg_pkg::ecc_reg__in_t hwif_in,
        output ecc_reg_pkg::ecc_reg__out_t hwif_out
    );

    //--------------------------------------------------------------------------
    // CPU Bus interface logic
    //--------------------------------------------------------------------------
    logic cpuif_req;
    logic cpuif_req_is_wr;
    logic [10:0] cpuif_addr;
    logic [31:0] cpuif_wr_data;
    logic cpuif_req_stall_wr;
    logic cpuif_req_stall_rd;

    logic cpuif_rd_ack;
    logic cpuif_rd_err;
    logic [31:0] cpuif_rd_data;

    logic cpuif_wr_ack;
    logic cpuif_wr_err;

    assign cpuif_req = s_cpuif_req;
    assign cpuif_req_is_wr = s_cpuif_req_is_wr;
    assign cpuif_addr = s_cpuif_addr;
    assign cpuif_wr_data = s_cpuif_wr_data;
    assign s_cpuif_req_stall_wr = cpuif_req_stall_wr;
    assign s_cpuif_req_stall_rd = cpuif_req_stall_rd;
    assign s_cpuif_rd_ack = cpuif_rd_ack;
    assign s_cpuif_rd_err = cpuif_rd_err;
    assign s_cpuif_rd_data = cpuif_rd_data;
    assign s_cpuif_wr_ack = cpuif_wr_ack;
    assign s_cpuif_wr_err = cpuif_wr_err;

    logic cpuif_req_masked;

    // Read & write latencies are balanced. Stalls not required
    assign cpuif_req_stall_rd = '0;
    assign cpuif_req_stall_wr = '0;
    assign cpuif_req_masked = cpuif_req;

    //--------------------------------------------------------------------------
    // Address Decode
    //--------------------------------------------------------------------------
    typedef struct {
        logic ecc_NAME[2];
        logic ecc_VERSION[2];
        logic ecc_CTRL;
        logic ecc_STATUS;
        logic ecc_SEED[12];
        logic ecc_MSG[12];
        logic ecc_PRIVKEY[12];
        logic ecc_PUBKEY_X[12];
        logic ecc_PUBKEY_Y[12];
        logic ecc_R[12];
        logic ecc_S[12];
        logic ecc_VERIFY_R[12];
        logic ecc_IV[12];
    } decoded_reg_strb_t;
    decoded_reg_strb_t decoded_reg_strb;
    logic decoded_req;
    logic decoded_req_is_wr;
    logic [31:0] decoded_wr_data;

    always_comb begin
        for(int i0=0; i0<2; i0++) begin
            decoded_reg_strb.ecc_NAME[i0] = cpuif_req_masked & (cpuif_addr == 'h0 + i0*'h4);
        end
        for(int i0=0; i0<2; i0++) begin
            decoded_reg_strb.ecc_VERSION[i0] = cpuif_req_masked & (cpuif_addr == 'h8 + i0*'h4);
        end
        decoded_reg_strb.ecc_CTRL = cpuif_req_masked & (cpuif_addr == 'h10);
        decoded_reg_strb.ecc_STATUS = cpuif_req_masked & (cpuif_addr == 'h18);
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_SEED[i0] = cpuif_req_masked & (cpuif_addr == 'h80 + i0*'h4);
        end
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_MSG[i0] = cpuif_req_masked & (cpuif_addr == 'h100 + i0*'h4);
        end
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_PRIVKEY[i0] = cpuif_req_masked & (cpuif_addr == 'h180 + i0*'h4);
        end
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_PUBKEY_X[i0] = cpuif_req_masked & (cpuif_addr == 'h200 + i0*'h4);
        end
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_PUBKEY_Y[i0] = cpuif_req_masked & (cpuif_addr == 'h280 + i0*'h4);
        end
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_R[i0] = cpuif_req_masked & (cpuif_addr == 'h300 + i0*'h4);
        end
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_S[i0] = cpuif_req_masked & (cpuif_addr == 'h380 + i0*'h4);
        end
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_VERIFY_R[i0] = cpuif_req_masked & (cpuif_addr == 'h400 + i0*'h4);
        end
        for(int i0=0; i0<12; i0++) begin
            decoded_reg_strb.ecc_IV[i0] = cpuif_req_masked & (cpuif_addr == 'h480 + i0*'h4);
        end
    end

    // Pass down signals to next stage
    assign decoded_req = cpuif_req_masked;
    assign decoded_req_is_wr = cpuif_req_is_wr;
    assign decoded_wr_data = cpuif_wr_data;

    // Writes are always granted with no error response
    assign cpuif_wr_ack = decoded_req & decoded_req_is_wr;
    assign cpuif_wr_err = '0;

    //--------------------------------------------------------------------------
    // Field logic
    //--------------------------------------------------------------------------
    typedef struct {
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } NAME;
        } ecc_NAME[2];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } VERSION;
        } ecc_VERSION[2];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } CTRL;
        } ecc_CTRL;
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } STATUS;
        } ecc_STATUS;
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } SEED;
        } ecc_SEED[12];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } MSG;
        } ecc_MSG[12];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } PRIVKEY;
        } ecc_PRIVKEY[12];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } PUBKEY_X;
        } ecc_PUBKEY_X[12];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } PUBKEY_Y;
        } ecc_PUBKEY_Y[12];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } R;
        } ecc_R[12];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } S;
        } ecc_S[12];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } VERIFY_R;
        } ecc_VERIFY_R[12];
        struct {
            struct {
                logic [31:0] next;
                logic load_next;
            } IV;
        } ecc_IV[12];
    } field_combo_t;
    field_combo_t field_combo;

    typedef struct {
        struct {
            struct {
                logic [31:0] value;
            } NAME;
        } ecc_NAME[2];
        struct {
            struct {
                logic [31:0] value;
            } VERSION;
        } ecc_VERSION[2];
        struct {
            struct {
                logic [31:0] value;
            } CTRL;
        } ecc_CTRL;
        struct {
            struct {
                logic [31:0] value;
            } STATUS;
        } ecc_STATUS;
        struct {
            struct {
                logic [31:0] value;
            } SEED;
        } ecc_SEED[12];
        struct {
            struct {
                logic [31:0] value;
            } MSG;
        } ecc_MSG[12];
        struct {
            struct {
                logic [31:0] value;
            } PRIVKEY;
        } ecc_PRIVKEY[12];
        struct {
            struct {
                logic [31:0] value;
            } PUBKEY_X;
        } ecc_PUBKEY_X[12];
        struct {
            struct {
                logic [31:0] value;
            } PUBKEY_Y;
        } ecc_PUBKEY_Y[12];
        struct {
            struct {
                logic [31:0] value;
            } R;
        } ecc_R[12];
        struct {
            struct {
                logic [31:0] value;
            } S;
        } ecc_S[12];
        struct {
            struct {
                logic [31:0] value;
            } VERIFY_R;
        } ecc_VERIFY_R[12];
        struct {
            struct {
                logic [31:0] value;
            } IV;
        } ecc_IV[12];
    } field_storage_t;
    field_storage_t field_storage;

    for(genvar i0=0; i0<2; i0++) begin
        // Field: ecc_reg.ecc_NAME[].NAME
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_NAME[i0].NAME.value;
            automatic logic load_next_c = '0;
            if(1) begin // HW Write
                next_c = hwif_in.ecc_NAME[i0].NAME.next;
                load_next_c = '1;
            end
            field_combo.ecc_NAME[i0].NAME.next = next_c;
            field_combo.ecc_NAME[i0].NAME.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_NAME[i0].NAME.load_next) begin
                field_storage.ecc_NAME[i0].NAME.value <= field_combo.ecc_NAME[i0].NAME.next;
            end
        end
        assign hwif_out.ecc_NAME[i0].NAME.value = field_storage.ecc_NAME[i0].NAME.value;
    end
    for(genvar i0=0; i0<2; i0++) begin
        // Field: ecc_reg.ecc_VERSION[].VERSION
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_VERSION[i0].VERSION.value;
            automatic logic load_next_c = '0;
            if(1) begin // HW Write
                next_c = hwif_in.ecc_VERSION[i0].VERSION.next;
                load_next_c = '1;
            end
            field_combo.ecc_VERSION[i0].VERSION.next = next_c;
            field_combo.ecc_VERSION[i0].VERSION.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_VERSION[i0].VERSION.load_next) begin
                field_storage.ecc_VERSION[i0].VERSION.value <= field_combo.ecc_VERSION[i0].VERSION.next;
            end
        end
        assign hwif_out.ecc_VERSION[i0].VERSION.value = field_storage.ecc_VERSION[i0].VERSION.value;
    end
    // Field: ecc_reg.ecc_CTRL.CTRL
    always_comb begin
        automatic logic [31:0] next_c = field_storage.ecc_CTRL.CTRL.value;
        automatic logic load_next_c = '0;
        if(decoded_reg_strb.ecc_CTRL && decoded_req_is_wr) begin // SW write
            next_c = decoded_wr_data[31:0];
            load_next_c = '1;
        end else if(1) begin // HW Write
            next_c = hwif_in.ecc_CTRL.CTRL.next;
            load_next_c = '1;
        end
        field_combo.ecc_CTRL.CTRL.next = next_c;
        field_combo.ecc_CTRL.CTRL.load_next = load_next_c;
    end
    always_ff @(posedge clk) begin
        if(field_combo.ecc_CTRL.CTRL.load_next) begin
            field_storage.ecc_CTRL.CTRL.value <= field_combo.ecc_CTRL.CTRL.next;
        end
    end
    assign hwif_out.ecc_CTRL.CTRL.value = field_storage.ecc_CTRL.CTRL.value;
    // Field: ecc_reg.ecc_STATUS.STATUS
    always_comb begin
        automatic logic [31:0] next_c = field_storage.ecc_STATUS.STATUS.value;
        automatic logic load_next_c = '0;
        if(1) begin // HW Write
            next_c = hwif_in.ecc_STATUS.STATUS.next;
            load_next_c = '1;
        end
        field_combo.ecc_STATUS.STATUS.next = next_c;
        field_combo.ecc_STATUS.STATUS.load_next = load_next_c;
    end
    always_ff @(posedge clk) begin
        if(field_combo.ecc_STATUS.STATUS.load_next) begin
            field_storage.ecc_STATUS.STATUS.value <= field_combo.ecc_STATUS.STATUS.next;
        end
    end
    assign hwif_out.ecc_STATUS.STATUS.value = field_storage.ecc_STATUS.STATUS.value;
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_SEED[].SEED
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_SEED[i0].SEED.value;
            automatic logic load_next_c = '0;
            if(decoded_reg_strb.ecc_SEED[i0] && decoded_req_is_wr) begin // SW write
                next_c = decoded_wr_data[31:0];
                load_next_c = '1;
            end else if(1) begin // HW Write
                next_c = hwif_in.ecc_SEED[i0].SEED.next;
                load_next_c = '1;
            end
            field_combo.ecc_SEED[i0].SEED.next = next_c;
            field_combo.ecc_SEED[i0].SEED.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_SEED[i0].SEED.load_next) begin
                field_storage.ecc_SEED[i0].SEED.value <= field_combo.ecc_SEED[i0].SEED.next;
            end
        end
        assign hwif_out.ecc_SEED[i0].SEED.value = field_storage.ecc_SEED[i0].SEED.value;
    end
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_MSG[].MSG
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_MSG[i0].MSG.value;
            automatic logic load_next_c = '0;
            if(decoded_reg_strb.ecc_MSG[i0] && decoded_req_is_wr) begin // SW write
                next_c = decoded_wr_data[31:0];
                load_next_c = '1;
            end
            field_combo.ecc_MSG[i0].MSG.next = next_c;
            field_combo.ecc_MSG[i0].MSG.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_MSG[i0].MSG.load_next) begin
                field_storage.ecc_MSG[i0].MSG.value <= field_combo.ecc_MSG[i0].MSG.next;
            end
        end
        assign hwif_out.ecc_MSG[i0].MSG.value = field_storage.ecc_MSG[i0].MSG.value;
    end
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_PRIVKEY[].PRIVKEY
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_PRIVKEY[i0].PRIVKEY.value;
            automatic logic load_next_c = '0;
            if(decoded_reg_strb.ecc_PRIVKEY[i0] && decoded_req_is_wr) begin // SW write
                next_c = decoded_wr_data[31:0];
                load_next_c = '1;
            end else if(1) begin // HW Write
                next_c = hwif_in.ecc_PRIVKEY[i0].PRIVKEY.next;
                load_next_c = '1;
            end
            field_combo.ecc_PRIVKEY[i0].PRIVKEY.next = next_c;
            field_combo.ecc_PRIVKEY[i0].PRIVKEY.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_PRIVKEY[i0].PRIVKEY.load_next) begin
                field_storage.ecc_PRIVKEY[i0].PRIVKEY.value <= field_combo.ecc_PRIVKEY[i0].PRIVKEY.next;
            end
        end
        assign hwif_out.ecc_PRIVKEY[i0].PRIVKEY.value = field_storage.ecc_PRIVKEY[i0].PRIVKEY.value;
    end
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_PUBKEY_X[].PUBKEY_X
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_PUBKEY_X[i0].PUBKEY_X.value;
            automatic logic load_next_c = '0;
            if(decoded_reg_strb.ecc_PUBKEY_X[i0] && decoded_req_is_wr) begin // SW write
                next_c = decoded_wr_data[31:0];
                load_next_c = '1;
            end else if(1) begin // HW Write
                next_c = hwif_in.ecc_PUBKEY_X[i0].PUBKEY_X.next;
                load_next_c = '1;
            end
            field_combo.ecc_PUBKEY_X[i0].PUBKEY_X.next = next_c;
            field_combo.ecc_PUBKEY_X[i0].PUBKEY_X.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_PUBKEY_X[i0].PUBKEY_X.load_next) begin
                field_storage.ecc_PUBKEY_X[i0].PUBKEY_X.value <= field_combo.ecc_PUBKEY_X[i0].PUBKEY_X.next;
            end
        end
        assign hwif_out.ecc_PUBKEY_X[i0].PUBKEY_X.value = field_storage.ecc_PUBKEY_X[i0].PUBKEY_X.value;
    end
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_PUBKEY_Y[].PUBKEY_Y
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_PUBKEY_Y[i0].PUBKEY_Y.value;
            automatic logic load_next_c = '0;
            if(decoded_reg_strb.ecc_PUBKEY_Y[i0] && decoded_req_is_wr) begin // SW write
                next_c = decoded_wr_data[31:0];
                load_next_c = '1;
            end else if(1) begin // HW Write
                next_c = hwif_in.ecc_PUBKEY_Y[i0].PUBKEY_Y.next;
                load_next_c = '1;
            end
            field_combo.ecc_PUBKEY_Y[i0].PUBKEY_Y.next = next_c;
            field_combo.ecc_PUBKEY_Y[i0].PUBKEY_Y.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_PUBKEY_Y[i0].PUBKEY_Y.load_next) begin
                field_storage.ecc_PUBKEY_Y[i0].PUBKEY_Y.value <= field_combo.ecc_PUBKEY_Y[i0].PUBKEY_Y.next;
            end
        end
        assign hwif_out.ecc_PUBKEY_Y[i0].PUBKEY_Y.value = field_storage.ecc_PUBKEY_Y[i0].PUBKEY_Y.value;
    end
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_R[].R
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_R[i0].R.value;
            automatic logic load_next_c = '0;
            if(decoded_reg_strb.ecc_R[i0] && decoded_req_is_wr) begin // SW write
                next_c = decoded_wr_data[31:0];
                load_next_c = '1;
            end else if(1) begin // HW Write
                next_c = hwif_in.ecc_R[i0].R.next;
                load_next_c = '1;
            end
            field_combo.ecc_R[i0].R.next = next_c;
            field_combo.ecc_R[i0].R.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_R[i0].R.load_next) begin
                field_storage.ecc_R[i0].R.value <= field_combo.ecc_R[i0].R.next;
            end
        end
        assign hwif_out.ecc_R[i0].R.value = field_storage.ecc_R[i0].R.value;
    end
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_S[].S
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_S[i0].S.value;
            automatic logic load_next_c = '0;
            if(decoded_reg_strb.ecc_S[i0] && decoded_req_is_wr) begin // SW write
                next_c = decoded_wr_data[31:0];
                load_next_c = '1;
            end else if(1) begin // HW Write
                next_c = hwif_in.ecc_S[i0].S.next;
                load_next_c = '1;
            end
            field_combo.ecc_S[i0].S.next = next_c;
            field_combo.ecc_S[i0].S.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_S[i0].S.load_next) begin
                field_storage.ecc_S[i0].S.value <= field_combo.ecc_S[i0].S.next;
            end
        end
        assign hwif_out.ecc_S[i0].S.value = field_storage.ecc_S[i0].S.value;
    end
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_VERIFY_R[].VERIFY_R
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_VERIFY_R[i0].VERIFY_R.value;
            automatic logic load_next_c = '0;
            if(1) begin // HW Write
                next_c = hwif_in.ecc_VERIFY_R[i0].VERIFY_R.next;
                load_next_c = '1;
            end
            field_combo.ecc_VERIFY_R[i0].VERIFY_R.next = next_c;
            field_combo.ecc_VERIFY_R[i0].VERIFY_R.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_VERIFY_R[i0].VERIFY_R.load_next) begin
                field_storage.ecc_VERIFY_R[i0].VERIFY_R.value <= field_combo.ecc_VERIFY_R[i0].VERIFY_R.next;
            end
        end
        assign hwif_out.ecc_VERIFY_R[i0].VERIFY_R.value = field_storage.ecc_VERIFY_R[i0].VERIFY_R.value;
    end
    for(genvar i0=0; i0<12; i0++) begin
        // Field: ecc_reg.ecc_IV[].IV
        always_comb begin
            automatic logic [31:0] next_c = field_storage.ecc_IV[i0].IV.value;
            automatic logic load_next_c = '0;
            if(decoded_reg_strb.ecc_IV[i0] && decoded_req_is_wr) begin // SW write
                next_c = decoded_wr_data[31:0];
                load_next_c = '1;
            end
            field_combo.ecc_IV[i0].IV.next = next_c;
            field_combo.ecc_IV[i0].IV.load_next = load_next_c;
        end
        always_ff @(posedge clk) begin
            if(field_combo.ecc_IV[i0].IV.load_next) begin
                field_storage.ecc_IV[i0].IV.value <= field_combo.ecc_IV[i0].IV.next;
            end
        end
        assign hwif_out.ecc_IV[i0].IV.value = field_storage.ecc_IV[i0].IV.value;
    end

    //--------------------------------------------------------------------------
    // Readback
    //--------------------------------------------------------------------------
    logic readback_err;
    logic readback_done;
    logic [31:0] readback_data;
    
    // Assign readback values to a flattened array
    logic [31:0] readback_array[114];
    for(genvar i0=0; i0<2; i0++) begin
        assign readback_array[i0*1 + 0][31:0] = (decoded_reg_strb.ecc_NAME[i0] && !decoded_req_is_wr) ? field_storage.ecc_NAME[i0].NAME.value : '0;
    end
    for(genvar i0=0; i0<2; i0++) begin
        assign readback_array[i0*1 + 2][31:0] = (decoded_reg_strb.ecc_VERSION[i0] && !decoded_req_is_wr) ? field_storage.ecc_VERSION[i0].VERSION.value : '0;
    end
    assign readback_array[4][31:0] = (decoded_reg_strb.ecc_CTRL && !decoded_req_is_wr) ? field_storage.ecc_CTRL.CTRL.value : '0;
    assign readback_array[5][31:0] = (decoded_reg_strb.ecc_STATUS && !decoded_req_is_wr) ? field_storage.ecc_STATUS.STATUS.value : '0;
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 6][31:0] = (decoded_reg_strb.ecc_SEED[i0] && !decoded_req_is_wr) ? field_storage.ecc_SEED[i0].SEED.value : '0;
    end
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 18][31:0] = (decoded_reg_strb.ecc_MSG[i0] && !decoded_req_is_wr) ? field_storage.ecc_MSG[i0].MSG.value : '0;
    end
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 30][31:0] = (decoded_reg_strb.ecc_PRIVKEY[i0] && !decoded_req_is_wr) ? field_storage.ecc_PRIVKEY[i0].PRIVKEY.value : '0;
    end
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 42][31:0] = (decoded_reg_strb.ecc_PUBKEY_X[i0] && !decoded_req_is_wr) ? field_storage.ecc_PUBKEY_X[i0].PUBKEY_X.value : '0;
    end
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 54][31:0] = (decoded_reg_strb.ecc_PUBKEY_Y[i0] && !decoded_req_is_wr) ? field_storage.ecc_PUBKEY_Y[i0].PUBKEY_Y.value : '0;
    end
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 66][31:0] = (decoded_reg_strb.ecc_R[i0] && !decoded_req_is_wr) ? field_storage.ecc_R[i0].R.value : '0;
    end
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 78][31:0] = (decoded_reg_strb.ecc_S[i0] && !decoded_req_is_wr) ? field_storage.ecc_S[i0].S.value : '0;
    end
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 90][31:0] = (decoded_reg_strb.ecc_VERIFY_R[i0] && !decoded_req_is_wr) ? field_storage.ecc_VERIFY_R[i0].VERIFY_R.value : '0;
    end
    for(genvar i0=0; i0<12; i0++) begin
        assign readback_array[i0*1 + 102][31:0] = (decoded_reg_strb.ecc_IV[i0] && !decoded_req_is_wr) ? field_storage.ecc_IV[i0].IV.value : '0;
    end


    // Reduce the array
    always_comb begin
        automatic logic [31:0] readback_data_var;
        readback_done = decoded_req & ~decoded_req_is_wr;
        readback_err = '0;
        readback_data_var = '0;
        for(int i=0; i<114; i++) readback_data_var |= readback_array[i];
        readback_data = readback_data_var;
    end


    assign cpuif_rd_ack = readback_done;
    assign cpuif_rd_data = readback_data;
    assign cpuif_rd_err = readback_err;


endmodule