//
// File: qvip_ahb_lite_slave_pkg.sv
//
// Generated from Mentor VIP Configurator (20220406)
// Generated using Mentor VIP Library ( 2022.2 : 04/20/2022:16:06 )
//
package qvip_ahb_lite_slave_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    import addr_map_pkg::*;
    
    import qvip_ahb_lite_slave_params_pkg::*;
    import mvc_pkg::*;
    import mgc_ahb_seq_pkg::*;
    import mgc_ahb_v2_0_pkg::*;
    
    `include "qvip_ahb_lite_slave_env_config.svh"
    `include "qvip_ahb_lite_slave_env.svh"
    `include "qvip_ahb_lite_slave_vseq_base.svh"
    `include "qvip_ahb_lite_slave_test_base.svh"
    `include "qvip_ahb_lite_slave_example_vseq.svh"
endpackage: qvip_ahb_lite_slave_pkg
