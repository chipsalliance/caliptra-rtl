// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef CALIPTRA_REG_DEFINES_HEADER
`define CALIPTRA_REG_DEFINES_HEADER


`define CLP_BASE_ADDR                                                                               (32'h0)
`define CLP_DOE_REG_BASE_ADDR                                                                       (32'h10000000)
`define CLP_DOE_REG_DOE_IV_0                                                                        (32'h10000000)
`define DOE_REG_DOE_IV_0                                                                            (32'h0)
`define CLP_DOE_REG_DOE_IV_1                                                                        (32'h10000004)
`define DOE_REG_DOE_IV_1                                                                            (32'h4)
`define CLP_DOE_REG_DOE_IV_2                                                                        (32'h10000008)
`define DOE_REG_DOE_IV_2                                                                            (32'h8)
`define CLP_DOE_REG_DOE_IV_3                                                                        (32'h1000000c)
`define DOE_REG_DOE_IV_3                                                                            (32'hc)
`define CLP_DOE_REG_DOE_CTRL                                                                        (32'h10000010)
`define DOE_REG_DOE_CTRL                                                                            (32'h10)
`define DOE_REG_DOE_CTRL_CMD_LOW                                                                    (0)
`define DOE_REG_DOE_CTRL_CMD_MASK                                                                   (32'h3)
`define DOE_REG_DOE_CTRL_DEST_LOW                                                                   (2)
`define DOE_REG_DOE_CTRL_DEST_MASK                                                                  (32'h1c)
`define CLP_DOE_REG_DOE_STATUS                                                                      (32'h10000014)
`define DOE_REG_DOE_STATUS                                                                          (32'h14)
`define DOE_REG_DOE_STATUS_READY_LOW                                                                (0)
`define DOE_REG_DOE_STATUS_READY_MASK                                                               (32'h1)
`define DOE_REG_DOE_STATUS_VALID_LOW                                                                (1)
`define DOE_REG_DOE_STATUS_VALID_MASK                                                               (32'h2)
`define CLP_DOE_REG_INTR_BLOCK_RF_START                                                             (32'h10000800)
`define CLP_DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10000800)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                      (32'h800)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                         (0)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                        (32'h1)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                         (1)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                        (32'h2)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10000804)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                       (32'h804)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                         (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                        (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                         (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                        (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                         (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                        (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                         (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                        (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10000808)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                       (32'h808)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                 (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                                (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1000080c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                   (32'h80c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10000810)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                   (32'h810)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10000814)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                 (32'h814)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                                  (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                                 (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                                  (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                                 (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                                  (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                                 (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                                  (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                                 (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10000818)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                 (32'h818)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                          (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                         (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1000081c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                     (32'h81c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                     (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                    (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                     (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                    (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                     (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                    (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                     (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                    (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10000820)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                     (32'h820)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                             (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                            (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                               (32'h10000900)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                   (32'h900)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                               (32'h10000904)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                   (32'h904)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                               (32'h10000908)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                   (32'h908)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                               (32'h1000090c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                   (32'h90c)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10000980)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                           (32'h980)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                          (32'h10000a00)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                              (32'ha00)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                          (32'h10000a04)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                              (32'ha04)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                          (32'h10000a08)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                              (32'ha08)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                          (32'h10000a0c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                              (32'ha0c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10000a10)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                      (32'ha10)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_ECC_REG_BASE_ADDR                                                                       (32'h10008000)
`define CLP_ECC_REG_ECC_NAME_0                                                                      (32'h10008000)
`define ECC_REG_ECC_NAME_0                                                                          (32'h0)
`define CLP_ECC_REG_ECC_NAME_1                                                                      (32'h10008004)
`define ECC_REG_ECC_NAME_1                                                                          (32'h4)
`define CLP_ECC_REG_ECC_VERSION_0                                                                   (32'h10008008)
`define ECC_REG_ECC_VERSION_0                                                                       (32'h8)
`define CLP_ECC_REG_ECC_VERSION_1                                                                   (32'h1000800c)
`define ECC_REG_ECC_VERSION_1                                                                       (32'hc)
`define CLP_ECC_REG_ECC_CTRL                                                                        (32'h10008010)
`define ECC_REG_ECC_CTRL                                                                            (32'h10)
`define ECC_REG_ECC_CTRL_CTRL_LOW                                                                   (0)
`define ECC_REG_ECC_CTRL_CTRL_MASK                                                                  (32'h3)
`define ECC_REG_ECC_CTRL_ZEROIZE_LOW                                                                (2)
`define ECC_REG_ECC_CTRL_ZEROIZE_MASK                                                               (32'h4)
`define CLP_ECC_REG_ECC_STATUS                                                                      (32'h10008018)
`define ECC_REG_ECC_STATUS                                                                          (32'h18)
`define ECC_REG_ECC_STATUS_READY_LOW                                                                (0)
`define ECC_REG_ECC_STATUS_READY_MASK                                                               (32'h1)
`define ECC_REG_ECC_STATUS_VALID_LOW                                                                (1)
`define ECC_REG_ECC_STATUS_VALID_MASK                                                               (32'h2)
`define CLP_ECC_REG_ECC_SCACONFIG                                                                   (32'h10008020)
`define ECC_REG_ECC_SCACONFIG                                                                       (32'h20)
`define ECC_REG_ECC_SCACONFIG_POINT_RND_EN_LOW                                                      (0)
`define ECC_REG_ECC_SCACONFIG_POINT_RND_EN_MASK                                                     (32'h1)
`define ECC_REG_ECC_SCACONFIG_MASK_SIGN_EN_LOW                                                      (1)
`define ECC_REG_ECC_SCACONFIG_MASK_SIGN_EN_MASK                                                     (32'h2)
`define ECC_REG_ECC_SCACONFIG_SCALAR_RND_EN_LOW                                                     (2)
`define ECC_REG_ECC_SCACONFIG_SCALAR_RND_EN_MASK                                                    (32'h4)
`define CLP_ECC_REG_ECC_SEED_0                                                                      (32'h10008080)
`define ECC_REG_ECC_SEED_0                                                                          (32'h80)
`define CLP_ECC_REG_ECC_SEED_1                                                                      (32'h10008084)
`define ECC_REG_ECC_SEED_1                                                                          (32'h84)
`define CLP_ECC_REG_ECC_SEED_2                                                                      (32'h10008088)
`define ECC_REG_ECC_SEED_2                                                                          (32'h88)
`define CLP_ECC_REG_ECC_SEED_3                                                                      (32'h1000808c)
`define ECC_REG_ECC_SEED_3                                                                          (32'h8c)
`define CLP_ECC_REG_ECC_SEED_4                                                                      (32'h10008090)
`define ECC_REG_ECC_SEED_4                                                                          (32'h90)
`define CLP_ECC_REG_ECC_SEED_5                                                                      (32'h10008094)
`define ECC_REG_ECC_SEED_5                                                                          (32'h94)
`define CLP_ECC_REG_ECC_SEED_6                                                                      (32'h10008098)
`define ECC_REG_ECC_SEED_6                                                                          (32'h98)
`define CLP_ECC_REG_ECC_SEED_7                                                                      (32'h1000809c)
`define ECC_REG_ECC_SEED_7                                                                          (32'h9c)
`define CLP_ECC_REG_ECC_SEED_8                                                                      (32'h100080a0)
`define ECC_REG_ECC_SEED_8                                                                          (32'ha0)
`define CLP_ECC_REG_ECC_SEED_9                                                                      (32'h100080a4)
`define ECC_REG_ECC_SEED_9                                                                          (32'ha4)
`define CLP_ECC_REG_ECC_SEED_10                                                                     (32'h100080a8)
`define ECC_REG_ECC_SEED_10                                                                         (32'ha8)
`define CLP_ECC_REG_ECC_SEED_11                                                                     (32'h100080ac)
`define ECC_REG_ECC_SEED_11                                                                         (32'hac)
`define CLP_ECC_REG_ECC_MSG_0                                                                       (32'h10008100)
`define ECC_REG_ECC_MSG_0                                                                           (32'h100)
`define CLP_ECC_REG_ECC_MSG_1                                                                       (32'h10008104)
`define ECC_REG_ECC_MSG_1                                                                           (32'h104)
`define CLP_ECC_REG_ECC_MSG_2                                                                       (32'h10008108)
`define ECC_REG_ECC_MSG_2                                                                           (32'h108)
`define CLP_ECC_REG_ECC_MSG_3                                                                       (32'h1000810c)
`define ECC_REG_ECC_MSG_3                                                                           (32'h10c)
`define CLP_ECC_REG_ECC_MSG_4                                                                       (32'h10008110)
`define ECC_REG_ECC_MSG_4                                                                           (32'h110)
`define CLP_ECC_REG_ECC_MSG_5                                                                       (32'h10008114)
`define ECC_REG_ECC_MSG_5                                                                           (32'h114)
`define CLP_ECC_REG_ECC_MSG_6                                                                       (32'h10008118)
`define ECC_REG_ECC_MSG_6                                                                           (32'h118)
`define CLP_ECC_REG_ECC_MSG_7                                                                       (32'h1000811c)
`define ECC_REG_ECC_MSG_7                                                                           (32'h11c)
`define CLP_ECC_REG_ECC_MSG_8                                                                       (32'h10008120)
`define ECC_REG_ECC_MSG_8                                                                           (32'h120)
`define CLP_ECC_REG_ECC_MSG_9                                                                       (32'h10008124)
`define ECC_REG_ECC_MSG_9                                                                           (32'h124)
`define CLP_ECC_REG_ECC_MSG_10                                                                      (32'h10008128)
`define ECC_REG_ECC_MSG_10                                                                          (32'h128)
`define CLP_ECC_REG_ECC_MSG_11                                                                      (32'h1000812c)
`define ECC_REG_ECC_MSG_11                                                                          (32'h12c)
`define CLP_ECC_REG_ECC_PRIVKEY_0                                                                   (32'h10008180)
`define ECC_REG_ECC_PRIVKEY_0                                                                       (32'h180)
`define CLP_ECC_REG_ECC_PRIVKEY_1                                                                   (32'h10008184)
`define ECC_REG_ECC_PRIVKEY_1                                                                       (32'h184)
`define CLP_ECC_REG_ECC_PRIVKEY_2                                                                   (32'h10008188)
`define ECC_REG_ECC_PRIVKEY_2                                                                       (32'h188)
`define CLP_ECC_REG_ECC_PRIVKEY_3                                                                   (32'h1000818c)
`define ECC_REG_ECC_PRIVKEY_3                                                                       (32'h18c)
`define CLP_ECC_REG_ECC_PRIVKEY_4                                                                   (32'h10008190)
`define ECC_REG_ECC_PRIVKEY_4                                                                       (32'h190)
`define CLP_ECC_REG_ECC_PRIVKEY_5                                                                   (32'h10008194)
`define ECC_REG_ECC_PRIVKEY_5                                                                       (32'h194)
`define CLP_ECC_REG_ECC_PRIVKEY_6                                                                   (32'h10008198)
`define ECC_REG_ECC_PRIVKEY_6                                                                       (32'h198)
`define CLP_ECC_REG_ECC_PRIVKEY_7                                                                   (32'h1000819c)
`define ECC_REG_ECC_PRIVKEY_7                                                                       (32'h19c)
`define CLP_ECC_REG_ECC_PRIVKEY_8                                                                   (32'h100081a0)
`define ECC_REG_ECC_PRIVKEY_8                                                                       (32'h1a0)
`define CLP_ECC_REG_ECC_PRIVKEY_9                                                                   (32'h100081a4)
`define ECC_REG_ECC_PRIVKEY_9                                                                       (32'h1a4)
`define CLP_ECC_REG_ECC_PRIVKEY_10                                                                  (32'h100081a8)
`define ECC_REG_ECC_PRIVKEY_10                                                                      (32'h1a8)
`define CLP_ECC_REG_ECC_PRIVKEY_11                                                                  (32'h100081ac)
`define ECC_REG_ECC_PRIVKEY_11                                                                      (32'h1ac)
`define CLP_ECC_REG_ECC_PUBKEY_X_0                                                                  (32'h10008200)
`define ECC_REG_ECC_PUBKEY_X_0                                                                      (32'h200)
`define CLP_ECC_REG_ECC_PUBKEY_X_1                                                                  (32'h10008204)
`define ECC_REG_ECC_PUBKEY_X_1                                                                      (32'h204)
`define CLP_ECC_REG_ECC_PUBKEY_X_2                                                                  (32'h10008208)
`define ECC_REG_ECC_PUBKEY_X_2                                                                      (32'h208)
`define CLP_ECC_REG_ECC_PUBKEY_X_3                                                                  (32'h1000820c)
`define ECC_REG_ECC_PUBKEY_X_3                                                                      (32'h20c)
`define CLP_ECC_REG_ECC_PUBKEY_X_4                                                                  (32'h10008210)
`define ECC_REG_ECC_PUBKEY_X_4                                                                      (32'h210)
`define CLP_ECC_REG_ECC_PUBKEY_X_5                                                                  (32'h10008214)
`define ECC_REG_ECC_PUBKEY_X_5                                                                      (32'h214)
`define CLP_ECC_REG_ECC_PUBKEY_X_6                                                                  (32'h10008218)
`define ECC_REG_ECC_PUBKEY_X_6                                                                      (32'h218)
`define CLP_ECC_REG_ECC_PUBKEY_X_7                                                                  (32'h1000821c)
`define ECC_REG_ECC_PUBKEY_X_7                                                                      (32'h21c)
`define CLP_ECC_REG_ECC_PUBKEY_X_8                                                                  (32'h10008220)
`define ECC_REG_ECC_PUBKEY_X_8                                                                      (32'h220)
`define CLP_ECC_REG_ECC_PUBKEY_X_9                                                                  (32'h10008224)
`define ECC_REG_ECC_PUBKEY_X_9                                                                      (32'h224)
`define CLP_ECC_REG_ECC_PUBKEY_X_10                                                                 (32'h10008228)
`define ECC_REG_ECC_PUBKEY_X_10                                                                     (32'h228)
`define CLP_ECC_REG_ECC_PUBKEY_X_11                                                                 (32'h1000822c)
`define ECC_REG_ECC_PUBKEY_X_11                                                                     (32'h22c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_0                                                                  (32'h10008280)
`define ECC_REG_ECC_PUBKEY_Y_0                                                                      (32'h280)
`define CLP_ECC_REG_ECC_PUBKEY_Y_1                                                                  (32'h10008284)
`define ECC_REG_ECC_PUBKEY_Y_1                                                                      (32'h284)
`define CLP_ECC_REG_ECC_PUBKEY_Y_2                                                                  (32'h10008288)
`define ECC_REG_ECC_PUBKEY_Y_2                                                                      (32'h288)
`define CLP_ECC_REG_ECC_PUBKEY_Y_3                                                                  (32'h1000828c)
`define ECC_REG_ECC_PUBKEY_Y_3                                                                      (32'h28c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_4                                                                  (32'h10008290)
`define ECC_REG_ECC_PUBKEY_Y_4                                                                      (32'h290)
`define CLP_ECC_REG_ECC_PUBKEY_Y_5                                                                  (32'h10008294)
`define ECC_REG_ECC_PUBKEY_Y_5                                                                      (32'h294)
`define CLP_ECC_REG_ECC_PUBKEY_Y_6                                                                  (32'h10008298)
`define ECC_REG_ECC_PUBKEY_Y_6                                                                      (32'h298)
`define CLP_ECC_REG_ECC_PUBKEY_Y_7                                                                  (32'h1000829c)
`define ECC_REG_ECC_PUBKEY_Y_7                                                                      (32'h29c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_8                                                                  (32'h100082a0)
`define ECC_REG_ECC_PUBKEY_Y_8                                                                      (32'h2a0)
`define CLP_ECC_REG_ECC_PUBKEY_Y_9                                                                  (32'h100082a4)
`define ECC_REG_ECC_PUBKEY_Y_9                                                                      (32'h2a4)
`define CLP_ECC_REG_ECC_PUBKEY_Y_10                                                                 (32'h100082a8)
`define ECC_REG_ECC_PUBKEY_Y_10                                                                     (32'h2a8)
`define CLP_ECC_REG_ECC_PUBKEY_Y_11                                                                 (32'h100082ac)
`define ECC_REG_ECC_PUBKEY_Y_11                                                                     (32'h2ac)
`define CLP_ECC_REG_ECC_SIGN_R_0                                                                    (32'h10008300)
`define ECC_REG_ECC_SIGN_R_0                                                                        (32'h300)
`define CLP_ECC_REG_ECC_SIGN_R_1                                                                    (32'h10008304)
`define ECC_REG_ECC_SIGN_R_1                                                                        (32'h304)
`define CLP_ECC_REG_ECC_SIGN_R_2                                                                    (32'h10008308)
`define ECC_REG_ECC_SIGN_R_2                                                                        (32'h308)
`define CLP_ECC_REG_ECC_SIGN_R_3                                                                    (32'h1000830c)
`define ECC_REG_ECC_SIGN_R_3                                                                        (32'h30c)
`define CLP_ECC_REG_ECC_SIGN_R_4                                                                    (32'h10008310)
`define ECC_REG_ECC_SIGN_R_4                                                                        (32'h310)
`define CLP_ECC_REG_ECC_SIGN_R_5                                                                    (32'h10008314)
`define ECC_REG_ECC_SIGN_R_5                                                                        (32'h314)
`define CLP_ECC_REG_ECC_SIGN_R_6                                                                    (32'h10008318)
`define ECC_REG_ECC_SIGN_R_6                                                                        (32'h318)
`define CLP_ECC_REG_ECC_SIGN_R_7                                                                    (32'h1000831c)
`define ECC_REG_ECC_SIGN_R_7                                                                        (32'h31c)
`define CLP_ECC_REG_ECC_SIGN_R_8                                                                    (32'h10008320)
`define ECC_REG_ECC_SIGN_R_8                                                                        (32'h320)
`define CLP_ECC_REG_ECC_SIGN_R_9                                                                    (32'h10008324)
`define ECC_REG_ECC_SIGN_R_9                                                                        (32'h324)
`define CLP_ECC_REG_ECC_SIGN_R_10                                                                   (32'h10008328)
`define ECC_REG_ECC_SIGN_R_10                                                                       (32'h328)
`define CLP_ECC_REG_ECC_SIGN_R_11                                                                   (32'h1000832c)
`define ECC_REG_ECC_SIGN_R_11                                                                       (32'h32c)
`define CLP_ECC_REG_ECC_SIGN_S_0                                                                    (32'h10008380)
`define ECC_REG_ECC_SIGN_S_0                                                                        (32'h380)
`define CLP_ECC_REG_ECC_SIGN_S_1                                                                    (32'h10008384)
`define ECC_REG_ECC_SIGN_S_1                                                                        (32'h384)
`define CLP_ECC_REG_ECC_SIGN_S_2                                                                    (32'h10008388)
`define ECC_REG_ECC_SIGN_S_2                                                                        (32'h388)
`define CLP_ECC_REG_ECC_SIGN_S_3                                                                    (32'h1000838c)
`define ECC_REG_ECC_SIGN_S_3                                                                        (32'h38c)
`define CLP_ECC_REG_ECC_SIGN_S_4                                                                    (32'h10008390)
`define ECC_REG_ECC_SIGN_S_4                                                                        (32'h390)
`define CLP_ECC_REG_ECC_SIGN_S_5                                                                    (32'h10008394)
`define ECC_REG_ECC_SIGN_S_5                                                                        (32'h394)
`define CLP_ECC_REG_ECC_SIGN_S_6                                                                    (32'h10008398)
`define ECC_REG_ECC_SIGN_S_6                                                                        (32'h398)
`define CLP_ECC_REG_ECC_SIGN_S_7                                                                    (32'h1000839c)
`define ECC_REG_ECC_SIGN_S_7                                                                        (32'h39c)
`define CLP_ECC_REG_ECC_SIGN_S_8                                                                    (32'h100083a0)
`define ECC_REG_ECC_SIGN_S_8                                                                        (32'h3a0)
`define CLP_ECC_REG_ECC_SIGN_S_9                                                                    (32'h100083a4)
`define ECC_REG_ECC_SIGN_S_9                                                                        (32'h3a4)
`define CLP_ECC_REG_ECC_SIGN_S_10                                                                   (32'h100083a8)
`define ECC_REG_ECC_SIGN_S_10                                                                       (32'h3a8)
`define CLP_ECC_REG_ECC_SIGN_S_11                                                                   (32'h100083ac)
`define ECC_REG_ECC_SIGN_S_11                                                                       (32'h3ac)
`define CLP_ECC_REG_ECC_VERIFY_R_0                                                                  (32'h10008400)
`define ECC_REG_ECC_VERIFY_R_0                                                                      (32'h400)
`define CLP_ECC_REG_ECC_VERIFY_R_1                                                                  (32'h10008404)
`define ECC_REG_ECC_VERIFY_R_1                                                                      (32'h404)
`define CLP_ECC_REG_ECC_VERIFY_R_2                                                                  (32'h10008408)
`define ECC_REG_ECC_VERIFY_R_2                                                                      (32'h408)
`define CLP_ECC_REG_ECC_VERIFY_R_3                                                                  (32'h1000840c)
`define ECC_REG_ECC_VERIFY_R_3                                                                      (32'h40c)
`define CLP_ECC_REG_ECC_VERIFY_R_4                                                                  (32'h10008410)
`define ECC_REG_ECC_VERIFY_R_4                                                                      (32'h410)
`define CLP_ECC_REG_ECC_VERIFY_R_5                                                                  (32'h10008414)
`define ECC_REG_ECC_VERIFY_R_5                                                                      (32'h414)
`define CLP_ECC_REG_ECC_VERIFY_R_6                                                                  (32'h10008418)
`define ECC_REG_ECC_VERIFY_R_6                                                                      (32'h418)
`define CLP_ECC_REG_ECC_VERIFY_R_7                                                                  (32'h1000841c)
`define ECC_REG_ECC_VERIFY_R_7                                                                      (32'h41c)
`define CLP_ECC_REG_ECC_VERIFY_R_8                                                                  (32'h10008420)
`define ECC_REG_ECC_VERIFY_R_8                                                                      (32'h420)
`define CLP_ECC_REG_ECC_VERIFY_R_9                                                                  (32'h10008424)
`define ECC_REG_ECC_VERIFY_R_9                                                                      (32'h424)
`define CLP_ECC_REG_ECC_VERIFY_R_10                                                                 (32'h10008428)
`define ECC_REG_ECC_VERIFY_R_10                                                                     (32'h428)
`define CLP_ECC_REG_ECC_VERIFY_R_11                                                                 (32'h1000842c)
`define ECC_REG_ECC_VERIFY_R_11                                                                     (32'h42c)
`define CLP_ECC_REG_ECC_IV_0                                                                        (32'h10008480)
`define ECC_REG_ECC_IV_0                                                                            (32'h480)
`define CLP_ECC_REG_ECC_IV_1                                                                        (32'h10008484)
`define ECC_REG_ECC_IV_1                                                                            (32'h484)
`define CLP_ECC_REG_ECC_IV_2                                                                        (32'h10008488)
`define ECC_REG_ECC_IV_2                                                                            (32'h488)
`define CLP_ECC_REG_ECC_IV_3                                                                        (32'h1000848c)
`define ECC_REG_ECC_IV_3                                                                            (32'h48c)
`define CLP_ECC_REG_ECC_IV_4                                                                        (32'h10008490)
`define ECC_REG_ECC_IV_4                                                                            (32'h490)
`define CLP_ECC_REG_ECC_IV_5                                                                        (32'h10008494)
`define ECC_REG_ECC_IV_5                                                                            (32'h494)
`define CLP_ECC_REG_ECC_IV_6                                                                        (32'h10008498)
`define ECC_REG_ECC_IV_6                                                                            (32'h498)
`define CLP_ECC_REG_ECC_IV_7                                                                        (32'h1000849c)
`define ECC_REG_ECC_IV_7                                                                            (32'h49c)
`define CLP_ECC_REG_ECC_IV_8                                                                        (32'h100084a0)
`define ECC_REG_ECC_IV_8                                                                            (32'h4a0)
`define CLP_ECC_REG_ECC_IV_9                                                                        (32'h100084a4)
`define ECC_REG_ECC_IV_9                                                                            (32'h4a4)
`define CLP_ECC_REG_ECC_IV_10                                                                       (32'h100084a8)
`define ECC_REG_ECC_IV_10                                                                           (32'h4a8)
`define CLP_ECC_REG_ECC_IV_11                                                                       (32'h100084ac)
`define ECC_REG_ECC_IV_11                                                                           (32'h4ac)
`define CLP_ECC_REG_ECC_KV_RD_PKEY_CTRL                                                             (32'h10008600)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL                                                                 (32'h600)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_EN_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_EN_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_ENTRY_LOW                                                  (1)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_ENTRY_MASK                                                 (32'he)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_ENTRY_IS_PCR_LOW                                                (4)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_ENTRY_IS_PCR_MASK                                               (32'h10)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_ENTRY_DATA_SIZE_LOW                                             (5)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_ENTRY_DATA_SIZE_MASK                                            (32'h3e0)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_RSVD_LOW                                                        (10)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_RSVD_MASK                                                       (32'h3ffffc00)
`define CLP_ECC_REG_ECC_KV_RD_PKEY_STATUS                                                           (32'h10008604)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS                                                               (32'h604)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_ECC_KV_RD_SEED_CTRL                                                             (32'h10008608)
`define ECC_REG_ECC_KV_RD_SEED_CTRL                                                                 (32'h608)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_EN_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_EN_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_ENTRY_LOW                                                  (1)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_ENTRY_MASK                                                 (32'he)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_ENTRY_IS_PCR_LOW                                                (4)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_ENTRY_IS_PCR_MASK                                               (32'h10)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_ENTRY_DATA_SIZE_LOW                                             (5)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_ENTRY_DATA_SIZE_MASK                                            (32'h3e0)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_RSVD_LOW                                                        (10)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_RSVD_MASK                                                       (32'h3ffffc00)
`define CLP_ECC_REG_ECC_KV_RD_SEED_STATUS                                                           (32'h1000860c)
`define ECC_REG_ECC_KV_RD_SEED_STATUS                                                               (32'h60c)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_ECC_KV_RD_MSG_CTRL                                                              (32'h10008610)
`define ECC_REG_ECC_KV_RD_MSG_CTRL                                                                  (32'h610)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_READ_EN_LOW                                                      (0)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_READ_EN_MASK                                                     (32'h1)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_READ_ENTRY_LOW                                                   (1)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_READ_ENTRY_MASK                                                  (32'he)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_ENTRY_IS_PCR_LOW                                                 (4)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_ENTRY_IS_PCR_MASK                                                (32'h10)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_ENTRY_DATA_SIZE_LOW                                              (5)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_ENTRY_DATA_SIZE_MASK                                             (32'h3e0)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_RSVD_LOW                                                         (10)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_RSVD_MASK                                                        (32'h3ffffc00)
`define CLP_ECC_REG_ECC_KV_RD_MSG_STATUS                                                            (32'h10008614)
`define ECC_REG_ECC_KV_RD_MSG_STATUS                                                                (32'h614)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_READY_LOW                                                      (0)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_READY_MASK                                                     (32'h1)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_VALID_LOW                                                      (1)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_VALID_MASK                                                     (32'h2)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_ERROR_LOW                                                      (2)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_ERROR_MASK                                                     (32'h3fc)
`define CLP_ECC_REG_ECC_KV_WR_PKEY_CTRL                                                             (32'h10008618)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL                                                                 (32'h618)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_EN_LOW                                                    (0)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_EN_MASK                                                   (32'h1)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_ENTRY_LOW                                                 (1)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_ENTRY_MASK                                                (32'he)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ENTRY_IS_PCR_LOW                                                (4)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ENTRY_IS_PCR_MASK                                               (32'h10)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_KEY_DEST_VALID_LOW                                         (5)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_KEY_DEST_VALID_MASK                                        (32'h20)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                       (6)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                      (32'h40)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_SHA_BLOCK_DEST_VALID_LOW                                        (7)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_SHA_BLOCK_DEST_VALID_MASK                                       (32'h80)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_PKEY_DEST_VALID_LOW                                         (8)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_PKEY_DEST_VALID_MASK                                        (32'h100)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_SEED_DEST_VALID_LOW                                         (9)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_SEED_DEST_VALID_MASK                                        (32'h200)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_MSG_DEST_VALID_LOW                                          (10)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_MSG_DEST_VALID_MASK                                         (32'h400)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_RSVD_LOW                                                        (11)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_RSVD_MASK                                                       (32'h3ffff800)
`define CLP_ECC_REG_ECC_KV_WR_PKEY_STATUS                                                           (32'h1000861c)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS                                                               (32'h61c)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_INTR_BLOCK_RF_START                                                             (32'h10008800)
`define CLP_ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10008800)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                      (32'h800)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                         (0)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                        (32'h1)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                         (1)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                        (32'h2)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10008804)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                       (32'h804)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_LOW                                 (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_MASK                                (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10008808)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                       (32'h808)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                 (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                                (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1000880c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                   (32'h80c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10008810)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                   (32'h810)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10008814)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                 (32'h814)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_LOW                          (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_MASK                         (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10008818)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                 (32'h818)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                          (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                         (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1000881c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                     (32'h81c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_LOW                             (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_MASK                            (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10008820)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                     (32'h820)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                             (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                            (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h10008900)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                           (32'h900)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10008980)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                           (32'h980)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'h10008a00)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                      (32'ha00)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10008a04)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                      (32'ha04)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_HMAC_REG_BASE_ADDR                                                                      (32'h10010000)
`define CLP_HMAC_REG_HMAC384_NAME_0                                                                 (32'h10010000)
`define HMAC_REG_HMAC384_NAME_0                                                                     (32'h0)
`define CLP_HMAC_REG_HMAC384_NAME_1                                                                 (32'h10010004)
`define HMAC_REG_HMAC384_NAME_1                                                                     (32'h4)
`define CLP_HMAC_REG_HMAC384_VERSION_0                                                              (32'h10010008)
`define HMAC_REG_HMAC384_VERSION_0                                                                  (32'h8)
`define CLP_HMAC_REG_HMAC384_VERSION_1                                                              (32'h1001000c)
`define HMAC_REG_HMAC384_VERSION_1                                                                  (32'hc)
`define CLP_HMAC_REG_HMAC384_CTRL                                                                   (32'h10010010)
`define HMAC_REG_HMAC384_CTRL                                                                       (32'h10)
`define HMAC_REG_HMAC384_CTRL_INIT_LOW                                                              (0)
`define HMAC_REG_HMAC384_CTRL_INIT_MASK                                                             (32'h1)
`define HMAC_REG_HMAC384_CTRL_NEXT_LOW                                                              (1)
`define HMAC_REG_HMAC384_CTRL_NEXT_MASK                                                             (32'h2)
`define HMAC_REG_HMAC384_CTRL_ZEROIZE_LOW                                                           (2)
`define HMAC_REG_HMAC384_CTRL_ZEROIZE_MASK                                                          (32'h4)
`define CLP_HMAC_REG_HMAC384_STATUS                                                                 (32'h10010018)
`define HMAC_REG_HMAC384_STATUS                                                                     (32'h18)
`define HMAC_REG_HMAC384_STATUS_READY_LOW                                                           (0)
`define HMAC_REG_HMAC384_STATUS_READY_MASK                                                          (32'h1)
`define HMAC_REG_HMAC384_STATUS_VALID_LOW                                                           (1)
`define HMAC_REG_HMAC384_STATUS_VALID_MASK                                                          (32'h2)
`define CLP_HMAC_REG_HMAC384_KEY_0                                                                  (32'h10010040)
`define HMAC_REG_HMAC384_KEY_0                                                                      (32'h40)
`define CLP_HMAC_REG_HMAC384_KEY_1                                                                  (32'h10010044)
`define HMAC_REG_HMAC384_KEY_1                                                                      (32'h44)
`define CLP_HMAC_REG_HMAC384_KEY_2                                                                  (32'h10010048)
`define HMAC_REG_HMAC384_KEY_2                                                                      (32'h48)
`define CLP_HMAC_REG_HMAC384_KEY_3                                                                  (32'h1001004c)
`define HMAC_REG_HMAC384_KEY_3                                                                      (32'h4c)
`define CLP_HMAC_REG_HMAC384_KEY_4                                                                  (32'h10010050)
`define HMAC_REG_HMAC384_KEY_4                                                                      (32'h50)
`define CLP_HMAC_REG_HMAC384_KEY_5                                                                  (32'h10010054)
`define HMAC_REG_HMAC384_KEY_5                                                                      (32'h54)
`define CLP_HMAC_REG_HMAC384_KEY_6                                                                  (32'h10010058)
`define HMAC_REG_HMAC384_KEY_6                                                                      (32'h58)
`define CLP_HMAC_REG_HMAC384_KEY_7                                                                  (32'h1001005c)
`define HMAC_REG_HMAC384_KEY_7                                                                      (32'h5c)
`define CLP_HMAC_REG_HMAC384_KEY_8                                                                  (32'h10010060)
`define HMAC_REG_HMAC384_KEY_8                                                                      (32'h60)
`define CLP_HMAC_REG_HMAC384_KEY_9                                                                  (32'h10010064)
`define HMAC_REG_HMAC384_KEY_9                                                                      (32'h64)
`define CLP_HMAC_REG_HMAC384_KEY_10                                                                 (32'h10010068)
`define HMAC_REG_HMAC384_KEY_10                                                                     (32'h68)
`define CLP_HMAC_REG_HMAC384_KEY_11                                                                 (32'h1001006c)
`define HMAC_REG_HMAC384_KEY_11                                                                     (32'h6c)
`define CLP_HMAC_REG_HMAC384_BLOCK_0                                                                (32'h10010080)
`define HMAC_REG_HMAC384_BLOCK_0                                                                    (32'h80)
`define CLP_HMAC_REG_HMAC384_BLOCK_1                                                                (32'h10010084)
`define HMAC_REG_HMAC384_BLOCK_1                                                                    (32'h84)
`define CLP_HMAC_REG_HMAC384_BLOCK_2                                                                (32'h10010088)
`define HMAC_REG_HMAC384_BLOCK_2                                                                    (32'h88)
`define CLP_HMAC_REG_HMAC384_BLOCK_3                                                                (32'h1001008c)
`define HMAC_REG_HMAC384_BLOCK_3                                                                    (32'h8c)
`define CLP_HMAC_REG_HMAC384_BLOCK_4                                                                (32'h10010090)
`define HMAC_REG_HMAC384_BLOCK_4                                                                    (32'h90)
`define CLP_HMAC_REG_HMAC384_BLOCK_5                                                                (32'h10010094)
`define HMAC_REG_HMAC384_BLOCK_5                                                                    (32'h94)
`define CLP_HMAC_REG_HMAC384_BLOCK_6                                                                (32'h10010098)
`define HMAC_REG_HMAC384_BLOCK_6                                                                    (32'h98)
`define CLP_HMAC_REG_HMAC384_BLOCK_7                                                                (32'h1001009c)
`define HMAC_REG_HMAC384_BLOCK_7                                                                    (32'h9c)
`define CLP_HMAC_REG_HMAC384_BLOCK_8                                                                (32'h100100a0)
`define HMAC_REG_HMAC384_BLOCK_8                                                                    (32'ha0)
`define CLP_HMAC_REG_HMAC384_BLOCK_9                                                                (32'h100100a4)
`define HMAC_REG_HMAC384_BLOCK_9                                                                    (32'ha4)
`define CLP_HMAC_REG_HMAC384_BLOCK_10                                                               (32'h100100a8)
`define HMAC_REG_HMAC384_BLOCK_10                                                                   (32'ha8)
`define CLP_HMAC_REG_HMAC384_BLOCK_11                                                               (32'h100100ac)
`define HMAC_REG_HMAC384_BLOCK_11                                                                   (32'hac)
`define CLP_HMAC_REG_HMAC384_BLOCK_12                                                               (32'h100100b0)
`define HMAC_REG_HMAC384_BLOCK_12                                                                   (32'hb0)
`define CLP_HMAC_REG_HMAC384_BLOCK_13                                                               (32'h100100b4)
`define HMAC_REG_HMAC384_BLOCK_13                                                                   (32'hb4)
`define CLP_HMAC_REG_HMAC384_BLOCK_14                                                               (32'h100100b8)
`define HMAC_REG_HMAC384_BLOCK_14                                                                   (32'hb8)
`define CLP_HMAC_REG_HMAC384_BLOCK_15                                                               (32'h100100bc)
`define HMAC_REG_HMAC384_BLOCK_15                                                                   (32'hbc)
`define CLP_HMAC_REG_HMAC384_BLOCK_16                                                               (32'h100100c0)
`define HMAC_REG_HMAC384_BLOCK_16                                                                   (32'hc0)
`define CLP_HMAC_REG_HMAC384_BLOCK_17                                                               (32'h100100c4)
`define HMAC_REG_HMAC384_BLOCK_17                                                                   (32'hc4)
`define CLP_HMAC_REG_HMAC384_BLOCK_18                                                               (32'h100100c8)
`define HMAC_REG_HMAC384_BLOCK_18                                                                   (32'hc8)
`define CLP_HMAC_REG_HMAC384_BLOCK_19                                                               (32'h100100cc)
`define HMAC_REG_HMAC384_BLOCK_19                                                                   (32'hcc)
`define CLP_HMAC_REG_HMAC384_BLOCK_20                                                               (32'h100100d0)
`define HMAC_REG_HMAC384_BLOCK_20                                                                   (32'hd0)
`define CLP_HMAC_REG_HMAC384_BLOCK_21                                                               (32'h100100d4)
`define HMAC_REG_HMAC384_BLOCK_21                                                                   (32'hd4)
`define CLP_HMAC_REG_HMAC384_BLOCK_22                                                               (32'h100100d8)
`define HMAC_REG_HMAC384_BLOCK_22                                                                   (32'hd8)
`define CLP_HMAC_REG_HMAC384_BLOCK_23                                                               (32'h100100dc)
`define HMAC_REG_HMAC384_BLOCK_23                                                                   (32'hdc)
`define CLP_HMAC_REG_HMAC384_BLOCK_24                                                               (32'h100100e0)
`define HMAC_REG_HMAC384_BLOCK_24                                                                   (32'he0)
`define CLP_HMAC_REG_HMAC384_BLOCK_25                                                               (32'h100100e4)
`define HMAC_REG_HMAC384_BLOCK_25                                                                   (32'he4)
`define CLP_HMAC_REG_HMAC384_BLOCK_26                                                               (32'h100100e8)
`define HMAC_REG_HMAC384_BLOCK_26                                                                   (32'he8)
`define CLP_HMAC_REG_HMAC384_BLOCK_27                                                               (32'h100100ec)
`define HMAC_REG_HMAC384_BLOCK_27                                                                   (32'hec)
`define CLP_HMAC_REG_HMAC384_BLOCK_28                                                               (32'h100100f0)
`define HMAC_REG_HMAC384_BLOCK_28                                                                   (32'hf0)
`define CLP_HMAC_REG_HMAC384_BLOCK_29                                                               (32'h100100f4)
`define HMAC_REG_HMAC384_BLOCK_29                                                                   (32'hf4)
`define CLP_HMAC_REG_HMAC384_BLOCK_30                                                               (32'h100100f8)
`define HMAC_REG_HMAC384_BLOCK_30                                                                   (32'hf8)
`define CLP_HMAC_REG_HMAC384_BLOCK_31                                                               (32'h100100fc)
`define HMAC_REG_HMAC384_BLOCK_31                                                                   (32'hfc)
`define CLP_HMAC_REG_HMAC384_TAG_0                                                                  (32'h10010100)
`define HMAC_REG_HMAC384_TAG_0                                                                      (32'h100)
`define CLP_HMAC_REG_HMAC384_TAG_1                                                                  (32'h10010104)
`define HMAC_REG_HMAC384_TAG_1                                                                      (32'h104)
`define CLP_HMAC_REG_HMAC384_TAG_2                                                                  (32'h10010108)
`define HMAC_REG_HMAC384_TAG_2                                                                      (32'h108)
`define CLP_HMAC_REG_HMAC384_TAG_3                                                                  (32'h1001010c)
`define HMAC_REG_HMAC384_TAG_3                                                                      (32'h10c)
`define CLP_HMAC_REG_HMAC384_TAG_4                                                                  (32'h10010110)
`define HMAC_REG_HMAC384_TAG_4                                                                      (32'h110)
`define CLP_HMAC_REG_HMAC384_TAG_5                                                                  (32'h10010114)
`define HMAC_REG_HMAC384_TAG_5                                                                      (32'h114)
`define CLP_HMAC_REG_HMAC384_TAG_6                                                                  (32'h10010118)
`define HMAC_REG_HMAC384_TAG_6                                                                      (32'h118)
`define CLP_HMAC_REG_HMAC384_TAG_7                                                                  (32'h1001011c)
`define HMAC_REG_HMAC384_TAG_7                                                                      (32'h11c)
`define CLP_HMAC_REG_HMAC384_TAG_8                                                                  (32'h10010120)
`define HMAC_REG_HMAC384_TAG_8                                                                      (32'h120)
`define CLP_HMAC_REG_HMAC384_TAG_9                                                                  (32'h10010124)
`define HMAC_REG_HMAC384_TAG_9                                                                      (32'h124)
`define CLP_HMAC_REG_HMAC384_TAG_10                                                                 (32'h10010128)
`define HMAC_REG_HMAC384_TAG_10                                                                     (32'h128)
`define CLP_HMAC_REG_HMAC384_TAG_11                                                                 (32'h1001012c)
`define HMAC_REG_HMAC384_TAG_11                                                                     (32'h12c)
`define CLP_HMAC_REG_HMAC384_KV_RD_KEY_CTRL                                                         (32'h10010600)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL                                                             (32'h600)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_READ_EN_LOW                                                 (0)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_READ_EN_MASK                                                (32'h1)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_READ_ENTRY_LOW                                              (1)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_READ_ENTRY_MASK                                             (32'he)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_ENTRY_IS_PCR_LOW                                            (4)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_ENTRY_IS_PCR_MASK                                           (32'h10)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_ENTRY_DATA_SIZE_LOW                                         (5)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_ENTRY_DATA_SIZE_MASK                                        (32'h3e0)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_RSVD_LOW                                                    (10)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_RSVD_MASK                                                   (32'h3ffffc00)
`define CLP_HMAC_REG_HMAC384_KV_RD_KEY_STATUS                                                       (32'h10010604)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS                                                           (32'h604)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_READY_LOW                                                 (0)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_READY_MASK                                                (32'h1)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_VALID_LOW                                                 (1)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_VALID_MASK                                                (32'h2)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_ERROR_LOW                                                 (2)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_ERROR_MASK                                                (32'h3fc)
`define CLP_HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL                                                       (32'h10010608)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL                                                           (32'h608)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_READ_EN_LOW                                               (0)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_READ_EN_MASK                                              (32'h1)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_READ_ENTRY_LOW                                            (1)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_READ_ENTRY_MASK                                           (32'he)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_ENTRY_IS_PCR_LOW                                          (4)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_ENTRY_IS_PCR_MASK                                         (32'h10)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_ENTRY_DATA_SIZE_LOW                                       (5)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_ENTRY_DATA_SIZE_MASK                                      (32'h3e0)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_RSVD_LOW                                                  (10)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_RSVD_MASK                                                 (32'h3ffffc00)
`define CLP_HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS                                                     (32'h1001060c)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS                                                         (32'h60c)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_READY_LOW                                               (0)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_READY_MASK                                              (32'h1)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_VALID_LOW                                               (1)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_VALID_MASK                                              (32'h2)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_ERROR_LOW                                               (2)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_ERROR_MASK                                              (32'h3fc)
`define CLP_HMAC_REG_HMAC384_KV_WR_CTRL                                                             (32'h10010610)
`define HMAC_REG_HMAC384_KV_WR_CTRL                                                                 (32'h610)
`define HMAC_REG_HMAC384_KV_WR_CTRL_WRITE_EN_LOW                                                    (0)
`define HMAC_REG_HMAC384_KV_WR_CTRL_WRITE_EN_MASK                                                   (32'h1)
`define HMAC_REG_HMAC384_KV_WR_CTRL_WRITE_ENTRY_LOW                                                 (1)
`define HMAC_REG_HMAC384_KV_WR_CTRL_WRITE_ENTRY_MASK                                                (32'he)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ENTRY_IS_PCR_LOW                                                (4)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ENTRY_IS_PCR_MASK                                               (32'h10)
`define HMAC_REG_HMAC384_KV_WR_CTRL_HMAC_KEY_DEST_VALID_LOW                                         (5)
`define HMAC_REG_HMAC384_KV_WR_CTRL_HMAC_KEY_DEST_VALID_MASK                                        (32'h20)
`define HMAC_REG_HMAC384_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                       (6)
`define HMAC_REG_HMAC384_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                      (32'h40)
`define HMAC_REG_HMAC384_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_LOW                                        (7)
`define HMAC_REG_HMAC384_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_MASK                                       (32'h80)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_PKEY_DEST_VALID_LOW                                         (8)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_PKEY_DEST_VALID_MASK                                        (32'h100)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_SEED_DEST_VALID_LOW                                         (9)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_SEED_DEST_VALID_MASK                                        (32'h200)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_MSG_DEST_VALID_LOW                                          (10)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_MSG_DEST_VALID_MASK                                         (32'h400)
`define HMAC_REG_HMAC384_KV_WR_CTRL_RSVD_LOW                                                        (11)
`define HMAC_REG_HMAC384_KV_WR_CTRL_RSVD_MASK                                                       (32'h3ffff800)
`define CLP_HMAC_REG_HMAC384_KV_WR_STATUS                                                           (32'h10010614)
`define HMAC_REG_HMAC384_KV_WR_STATUS                                                               (32'h614)
`define HMAC_REG_HMAC384_KV_WR_STATUS_READY_LOW                                                     (0)
`define HMAC_REG_HMAC384_KV_WR_STATUS_READY_MASK                                                    (32'h1)
`define HMAC_REG_HMAC384_KV_WR_STATUS_VALID_LOW                                                     (1)
`define HMAC_REG_HMAC384_KV_WR_STATUS_VALID_MASK                                                    (32'h2)
`define HMAC_REG_HMAC384_KV_WR_STATUS_ERROR_LOW                                                     (2)
`define HMAC_REG_HMAC384_KV_WR_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_HMAC_REG_INTR_BLOCK_RF_START                                                            (32'h10010800)
`define CLP_HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                 (32'h10010800)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                     (32'h800)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                        (0)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                       (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                        (1)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                       (32'h2)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                  (32'h10010804)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                      (32'h804)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                        (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                       (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                        (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                       (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                        (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                       (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                        (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                       (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                  (32'h10010808)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                      (32'h808)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                               (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                              (32'h1001080c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                  (32'h80c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                      (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                     (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                              (32'h10010810)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                  (32'h810)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                      (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                     (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                            (32'h10010814)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                (32'h814)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                                 (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                                (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                                 (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                                (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                                 (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                                (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                                 (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                                (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                            (32'h10010818)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                (32'h818)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                         (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                        (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                (32'h1001081c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                    (32'h81c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                    (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                   (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                    (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                   (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                    (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                   (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                    (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                   (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                (32'h10010820)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                    (32'h820)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                            (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                           (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                              (32'h10010900)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                  (32'h900)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                              (32'h10010904)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                  (32'h904)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                              (32'h10010908)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                  (32'h908)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                              (32'h1001090c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                  (32'h90c)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                      (32'h10010980)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                          (32'h980)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                         (32'h10010a00)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                             (32'ha00)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                         (32'h10010a04)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                             (32'ha04)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                         (32'h10010a08)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                             (32'ha08)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                         (32'h10010a0c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                             (32'ha0c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                 (32'h10010a10)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                     (32'ha10)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                           (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                          (32'h1)
`define CLP_KV_REG_BASE_ADDR                                                                        (32'h10018000)
`define CLP_KV_REG_PCR_CTRL_0                                                                       (32'h10018000)
`define KV_REG_PCR_CTRL_0                                                                           (32'h0)
`define KV_REG_PCR_CTRL_0_LOCK_WR_LOW                                                               (0)
`define KV_REG_PCR_CTRL_0_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_PCR_CTRL_0_LOCK_USE_LOW                                                              (1)
`define KV_REG_PCR_CTRL_0_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_PCR_CTRL_0_CLEAR_LOW                                                                 (2)
`define KV_REG_PCR_CTRL_0_CLEAR_MASK                                                                (32'h4)
`define KV_REG_PCR_CTRL_0_RSVD0_LOW                                                                 (3)
`define KV_REG_PCR_CTRL_0_RSVD0_MASK                                                                (32'h8)
`define KV_REG_PCR_CTRL_0_RSVD1_LOW                                                                 (4)
`define KV_REG_PCR_CTRL_0_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_PCR_CTRL_0_DEST_VALID_LOW                                                            (8)
`define KV_REG_PCR_CTRL_0_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_PCR_CTRL_0_RSVD_LOW                                                                  (14)
`define KV_REG_PCR_CTRL_0_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_PCR_CTRL_1                                                                       (32'h10018004)
`define KV_REG_PCR_CTRL_1                                                                           (32'h4)
`define KV_REG_PCR_CTRL_1_LOCK_WR_LOW                                                               (0)
`define KV_REG_PCR_CTRL_1_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_PCR_CTRL_1_LOCK_USE_LOW                                                              (1)
`define KV_REG_PCR_CTRL_1_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_PCR_CTRL_1_CLEAR_LOW                                                                 (2)
`define KV_REG_PCR_CTRL_1_CLEAR_MASK                                                                (32'h4)
`define KV_REG_PCR_CTRL_1_RSVD0_LOW                                                                 (3)
`define KV_REG_PCR_CTRL_1_RSVD0_MASK                                                                (32'h8)
`define KV_REG_PCR_CTRL_1_RSVD1_LOW                                                                 (4)
`define KV_REG_PCR_CTRL_1_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_PCR_CTRL_1_DEST_VALID_LOW                                                            (8)
`define KV_REG_PCR_CTRL_1_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_PCR_CTRL_1_RSVD_LOW                                                                  (14)
`define KV_REG_PCR_CTRL_1_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_PCR_CTRL_2                                                                       (32'h10018008)
`define KV_REG_PCR_CTRL_2                                                                           (32'h8)
`define KV_REG_PCR_CTRL_2_LOCK_WR_LOW                                                               (0)
`define KV_REG_PCR_CTRL_2_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_PCR_CTRL_2_LOCK_USE_LOW                                                              (1)
`define KV_REG_PCR_CTRL_2_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_PCR_CTRL_2_CLEAR_LOW                                                                 (2)
`define KV_REG_PCR_CTRL_2_CLEAR_MASK                                                                (32'h4)
`define KV_REG_PCR_CTRL_2_RSVD0_LOW                                                                 (3)
`define KV_REG_PCR_CTRL_2_RSVD0_MASK                                                                (32'h8)
`define KV_REG_PCR_CTRL_2_RSVD1_LOW                                                                 (4)
`define KV_REG_PCR_CTRL_2_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_PCR_CTRL_2_DEST_VALID_LOW                                                            (8)
`define KV_REG_PCR_CTRL_2_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_PCR_CTRL_2_RSVD_LOW                                                                  (14)
`define KV_REG_PCR_CTRL_2_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_PCR_CTRL_3                                                                       (32'h1001800c)
`define KV_REG_PCR_CTRL_3                                                                           (32'hc)
`define KV_REG_PCR_CTRL_3_LOCK_WR_LOW                                                               (0)
`define KV_REG_PCR_CTRL_3_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_PCR_CTRL_3_LOCK_USE_LOW                                                              (1)
`define KV_REG_PCR_CTRL_3_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_PCR_CTRL_3_CLEAR_LOW                                                                 (2)
`define KV_REG_PCR_CTRL_3_CLEAR_MASK                                                                (32'h4)
`define KV_REG_PCR_CTRL_3_RSVD0_LOW                                                                 (3)
`define KV_REG_PCR_CTRL_3_RSVD0_MASK                                                                (32'h8)
`define KV_REG_PCR_CTRL_3_RSVD1_LOW                                                                 (4)
`define KV_REG_PCR_CTRL_3_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_PCR_CTRL_3_DEST_VALID_LOW                                                            (8)
`define KV_REG_PCR_CTRL_3_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_PCR_CTRL_3_RSVD_LOW                                                                  (14)
`define KV_REG_PCR_CTRL_3_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_PCR_CTRL_4                                                                       (32'h10018010)
`define KV_REG_PCR_CTRL_4                                                                           (32'h10)
`define KV_REG_PCR_CTRL_4_LOCK_WR_LOW                                                               (0)
`define KV_REG_PCR_CTRL_4_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_PCR_CTRL_4_LOCK_USE_LOW                                                              (1)
`define KV_REG_PCR_CTRL_4_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_PCR_CTRL_4_CLEAR_LOW                                                                 (2)
`define KV_REG_PCR_CTRL_4_CLEAR_MASK                                                                (32'h4)
`define KV_REG_PCR_CTRL_4_RSVD0_LOW                                                                 (3)
`define KV_REG_PCR_CTRL_4_RSVD0_MASK                                                                (32'h8)
`define KV_REG_PCR_CTRL_4_RSVD1_LOW                                                                 (4)
`define KV_REG_PCR_CTRL_4_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_PCR_CTRL_4_DEST_VALID_LOW                                                            (8)
`define KV_REG_PCR_CTRL_4_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_PCR_CTRL_4_RSVD_LOW                                                                  (14)
`define KV_REG_PCR_CTRL_4_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_PCR_CTRL_5                                                                       (32'h10018014)
`define KV_REG_PCR_CTRL_5                                                                           (32'h14)
`define KV_REG_PCR_CTRL_5_LOCK_WR_LOW                                                               (0)
`define KV_REG_PCR_CTRL_5_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_PCR_CTRL_5_LOCK_USE_LOW                                                              (1)
`define KV_REG_PCR_CTRL_5_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_PCR_CTRL_5_CLEAR_LOW                                                                 (2)
`define KV_REG_PCR_CTRL_5_CLEAR_MASK                                                                (32'h4)
`define KV_REG_PCR_CTRL_5_RSVD0_LOW                                                                 (3)
`define KV_REG_PCR_CTRL_5_RSVD0_MASK                                                                (32'h8)
`define KV_REG_PCR_CTRL_5_RSVD1_LOW                                                                 (4)
`define KV_REG_PCR_CTRL_5_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_PCR_CTRL_5_DEST_VALID_LOW                                                            (8)
`define KV_REG_PCR_CTRL_5_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_PCR_CTRL_5_RSVD_LOW                                                                  (14)
`define KV_REG_PCR_CTRL_5_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_PCR_CTRL_6                                                                       (32'h10018018)
`define KV_REG_PCR_CTRL_6                                                                           (32'h18)
`define KV_REG_PCR_CTRL_6_LOCK_WR_LOW                                                               (0)
`define KV_REG_PCR_CTRL_6_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_PCR_CTRL_6_LOCK_USE_LOW                                                              (1)
`define KV_REG_PCR_CTRL_6_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_PCR_CTRL_6_CLEAR_LOW                                                                 (2)
`define KV_REG_PCR_CTRL_6_CLEAR_MASK                                                                (32'h4)
`define KV_REG_PCR_CTRL_6_RSVD0_LOW                                                                 (3)
`define KV_REG_PCR_CTRL_6_RSVD0_MASK                                                                (32'h8)
`define KV_REG_PCR_CTRL_6_RSVD1_LOW                                                                 (4)
`define KV_REG_PCR_CTRL_6_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_PCR_CTRL_6_DEST_VALID_LOW                                                            (8)
`define KV_REG_PCR_CTRL_6_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_PCR_CTRL_6_RSVD_LOW                                                                  (14)
`define KV_REG_PCR_CTRL_6_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_PCR_CTRL_7                                                                       (32'h1001801c)
`define KV_REG_PCR_CTRL_7                                                                           (32'h1c)
`define KV_REG_PCR_CTRL_7_LOCK_WR_LOW                                                               (0)
`define KV_REG_PCR_CTRL_7_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_PCR_CTRL_7_LOCK_USE_LOW                                                              (1)
`define KV_REG_PCR_CTRL_7_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_PCR_CTRL_7_CLEAR_LOW                                                                 (2)
`define KV_REG_PCR_CTRL_7_CLEAR_MASK                                                                (32'h4)
`define KV_REG_PCR_CTRL_7_RSVD0_LOW                                                                 (3)
`define KV_REG_PCR_CTRL_7_RSVD0_MASK                                                                (32'h8)
`define KV_REG_PCR_CTRL_7_RSVD1_LOW                                                                 (4)
`define KV_REG_PCR_CTRL_7_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_PCR_CTRL_7_DEST_VALID_LOW                                                            (8)
`define KV_REG_PCR_CTRL_7_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_PCR_CTRL_7_RSVD_LOW                                                                  (14)
`define KV_REG_PCR_CTRL_7_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_PCR_ENTRY_0_0                                                                    (32'h10018200)
`define KV_REG_PCR_ENTRY_0_0                                                                        (32'h200)
`define CLP_KV_REG_PCR_ENTRY_0_1                                                                    (32'h10018204)
`define KV_REG_PCR_ENTRY_0_1                                                                        (32'h204)
`define CLP_KV_REG_PCR_ENTRY_0_2                                                                    (32'h10018208)
`define KV_REG_PCR_ENTRY_0_2                                                                        (32'h208)
`define CLP_KV_REG_PCR_ENTRY_0_3                                                                    (32'h1001820c)
`define KV_REG_PCR_ENTRY_0_3                                                                        (32'h20c)
`define CLP_KV_REG_PCR_ENTRY_0_4                                                                    (32'h10018210)
`define KV_REG_PCR_ENTRY_0_4                                                                        (32'h210)
`define CLP_KV_REG_PCR_ENTRY_0_5                                                                    (32'h10018214)
`define KV_REG_PCR_ENTRY_0_5                                                                        (32'h214)
`define CLP_KV_REG_PCR_ENTRY_0_6                                                                    (32'h10018218)
`define KV_REG_PCR_ENTRY_0_6                                                                        (32'h218)
`define CLP_KV_REG_PCR_ENTRY_0_7                                                                    (32'h1001821c)
`define KV_REG_PCR_ENTRY_0_7                                                                        (32'h21c)
`define CLP_KV_REG_PCR_ENTRY_0_8                                                                    (32'h10018220)
`define KV_REG_PCR_ENTRY_0_8                                                                        (32'h220)
`define CLP_KV_REG_PCR_ENTRY_0_9                                                                    (32'h10018224)
`define KV_REG_PCR_ENTRY_0_9                                                                        (32'h224)
`define CLP_KV_REG_PCR_ENTRY_0_10                                                                   (32'h10018228)
`define KV_REG_PCR_ENTRY_0_10                                                                       (32'h228)
`define CLP_KV_REG_PCR_ENTRY_0_11                                                                   (32'h1001822c)
`define KV_REG_PCR_ENTRY_0_11                                                                       (32'h22c)
`define CLP_KV_REG_PCR_ENTRY_0_12                                                                   (32'h10018230)
`define KV_REG_PCR_ENTRY_0_12                                                                       (32'h230)
`define CLP_KV_REG_PCR_ENTRY_0_13                                                                   (32'h10018234)
`define KV_REG_PCR_ENTRY_0_13                                                                       (32'h234)
`define CLP_KV_REG_PCR_ENTRY_0_14                                                                   (32'h10018238)
`define KV_REG_PCR_ENTRY_0_14                                                                       (32'h238)
`define CLP_KV_REG_PCR_ENTRY_0_15                                                                   (32'h1001823c)
`define KV_REG_PCR_ENTRY_0_15                                                                       (32'h23c)
`define CLP_KV_REG_PCR_ENTRY_1_0                                                                    (32'h10018240)
`define KV_REG_PCR_ENTRY_1_0                                                                        (32'h240)
`define CLP_KV_REG_PCR_ENTRY_1_1                                                                    (32'h10018244)
`define KV_REG_PCR_ENTRY_1_1                                                                        (32'h244)
`define CLP_KV_REG_PCR_ENTRY_1_2                                                                    (32'h10018248)
`define KV_REG_PCR_ENTRY_1_2                                                                        (32'h248)
`define CLP_KV_REG_PCR_ENTRY_1_3                                                                    (32'h1001824c)
`define KV_REG_PCR_ENTRY_1_3                                                                        (32'h24c)
`define CLP_KV_REG_PCR_ENTRY_1_4                                                                    (32'h10018250)
`define KV_REG_PCR_ENTRY_1_4                                                                        (32'h250)
`define CLP_KV_REG_PCR_ENTRY_1_5                                                                    (32'h10018254)
`define KV_REG_PCR_ENTRY_1_5                                                                        (32'h254)
`define CLP_KV_REG_PCR_ENTRY_1_6                                                                    (32'h10018258)
`define KV_REG_PCR_ENTRY_1_6                                                                        (32'h258)
`define CLP_KV_REG_PCR_ENTRY_1_7                                                                    (32'h1001825c)
`define KV_REG_PCR_ENTRY_1_7                                                                        (32'h25c)
`define CLP_KV_REG_PCR_ENTRY_1_8                                                                    (32'h10018260)
`define KV_REG_PCR_ENTRY_1_8                                                                        (32'h260)
`define CLP_KV_REG_PCR_ENTRY_1_9                                                                    (32'h10018264)
`define KV_REG_PCR_ENTRY_1_9                                                                        (32'h264)
`define CLP_KV_REG_PCR_ENTRY_1_10                                                                   (32'h10018268)
`define KV_REG_PCR_ENTRY_1_10                                                                       (32'h268)
`define CLP_KV_REG_PCR_ENTRY_1_11                                                                   (32'h1001826c)
`define KV_REG_PCR_ENTRY_1_11                                                                       (32'h26c)
`define CLP_KV_REG_PCR_ENTRY_1_12                                                                   (32'h10018270)
`define KV_REG_PCR_ENTRY_1_12                                                                       (32'h270)
`define CLP_KV_REG_PCR_ENTRY_1_13                                                                   (32'h10018274)
`define KV_REG_PCR_ENTRY_1_13                                                                       (32'h274)
`define CLP_KV_REG_PCR_ENTRY_1_14                                                                   (32'h10018278)
`define KV_REG_PCR_ENTRY_1_14                                                                       (32'h278)
`define CLP_KV_REG_PCR_ENTRY_1_15                                                                   (32'h1001827c)
`define KV_REG_PCR_ENTRY_1_15                                                                       (32'h27c)
`define CLP_KV_REG_PCR_ENTRY_2_0                                                                    (32'h10018280)
`define KV_REG_PCR_ENTRY_2_0                                                                        (32'h280)
`define CLP_KV_REG_PCR_ENTRY_2_1                                                                    (32'h10018284)
`define KV_REG_PCR_ENTRY_2_1                                                                        (32'h284)
`define CLP_KV_REG_PCR_ENTRY_2_2                                                                    (32'h10018288)
`define KV_REG_PCR_ENTRY_2_2                                                                        (32'h288)
`define CLP_KV_REG_PCR_ENTRY_2_3                                                                    (32'h1001828c)
`define KV_REG_PCR_ENTRY_2_3                                                                        (32'h28c)
`define CLP_KV_REG_PCR_ENTRY_2_4                                                                    (32'h10018290)
`define KV_REG_PCR_ENTRY_2_4                                                                        (32'h290)
`define CLP_KV_REG_PCR_ENTRY_2_5                                                                    (32'h10018294)
`define KV_REG_PCR_ENTRY_2_5                                                                        (32'h294)
`define CLP_KV_REG_PCR_ENTRY_2_6                                                                    (32'h10018298)
`define KV_REG_PCR_ENTRY_2_6                                                                        (32'h298)
`define CLP_KV_REG_PCR_ENTRY_2_7                                                                    (32'h1001829c)
`define KV_REG_PCR_ENTRY_2_7                                                                        (32'h29c)
`define CLP_KV_REG_PCR_ENTRY_2_8                                                                    (32'h100182a0)
`define KV_REG_PCR_ENTRY_2_8                                                                        (32'h2a0)
`define CLP_KV_REG_PCR_ENTRY_2_9                                                                    (32'h100182a4)
`define KV_REG_PCR_ENTRY_2_9                                                                        (32'h2a4)
`define CLP_KV_REG_PCR_ENTRY_2_10                                                                   (32'h100182a8)
`define KV_REG_PCR_ENTRY_2_10                                                                       (32'h2a8)
`define CLP_KV_REG_PCR_ENTRY_2_11                                                                   (32'h100182ac)
`define KV_REG_PCR_ENTRY_2_11                                                                       (32'h2ac)
`define CLP_KV_REG_PCR_ENTRY_2_12                                                                   (32'h100182b0)
`define KV_REG_PCR_ENTRY_2_12                                                                       (32'h2b0)
`define CLP_KV_REG_PCR_ENTRY_2_13                                                                   (32'h100182b4)
`define KV_REG_PCR_ENTRY_2_13                                                                       (32'h2b4)
`define CLP_KV_REG_PCR_ENTRY_2_14                                                                   (32'h100182b8)
`define KV_REG_PCR_ENTRY_2_14                                                                       (32'h2b8)
`define CLP_KV_REG_PCR_ENTRY_2_15                                                                   (32'h100182bc)
`define KV_REG_PCR_ENTRY_2_15                                                                       (32'h2bc)
`define CLP_KV_REG_PCR_ENTRY_3_0                                                                    (32'h100182c0)
`define KV_REG_PCR_ENTRY_3_0                                                                        (32'h2c0)
`define CLP_KV_REG_PCR_ENTRY_3_1                                                                    (32'h100182c4)
`define KV_REG_PCR_ENTRY_3_1                                                                        (32'h2c4)
`define CLP_KV_REG_PCR_ENTRY_3_2                                                                    (32'h100182c8)
`define KV_REG_PCR_ENTRY_3_2                                                                        (32'h2c8)
`define CLP_KV_REG_PCR_ENTRY_3_3                                                                    (32'h100182cc)
`define KV_REG_PCR_ENTRY_3_3                                                                        (32'h2cc)
`define CLP_KV_REG_PCR_ENTRY_3_4                                                                    (32'h100182d0)
`define KV_REG_PCR_ENTRY_3_4                                                                        (32'h2d0)
`define CLP_KV_REG_PCR_ENTRY_3_5                                                                    (32'h100182d4)
`define KV_REG_PCR_ENTRY_3_5                                                                        (32'h2d4)
`define CLP_KV_REG_PCR_ENTRY_3_6                                                                    (32'h100182d8)
`define KV_REG_PCR_ENTRY_3_6                                                                        (32'h2d8)
`define CLP_KV_REG_PCR_ENTRY_3_7                                                                    (32'h100182dc)
`define KV_REG_PCR_ENTRY_3_7                                                                        (32'h2dc)
`define CLP_KV_REG_PCR_ENTRY_3_8                                                                    (32'h100182e0)
`define KV_REG_PCR_ENTRY_3_8                                                                        (32'h2e0)
`define CLP_KV_REG_PCR_ENTRY_3_9                                                                    (32'h100182e4)
`define KV_REG_PCR_ENTRY_3_9                                                                        (32'h2e4)
`define CLP_KV_REG_PCR_ENTRY_3_10                                                                   (32'h100182e8)
`define KV_REG_PCR_ENTRY_3_10                                                                       (32'h2e8)
`define CLP_KV_REG_PCR_ENTRY_3_11                                                                   (32'h100182ec)
`define KV_REG_PCR_ENTRY_3_11                                                                       (32'h2ec)
`define CLP_KV_REG_PCR_ENTRY_3_12                                                                   (32'h100182f0)
`define KV_REG_PCR_ENTRY_3_12                                                                       (32'h2f0)
`define CLP_KV_REG_PCR_ENTRY_3_13                                                                   (32'h100182f4)
`define KV_REG_PCR_ENTRY_3_13                                                                       (32'h2f4)
`define CLP_KV_REG_PCR_ENTRY_3_14                                                                   (32'h100182f8)
`define KV_REG_PCR_ENTRY_3_14                                                                       (32'h2f8)
`define CLP_KV_REG_PCR_ENTRY_3_15                                                                   (32'h100182fc)
`define KV_REG_PCR_ENTRY_3_15                                                                       (32'h2fc)
`define CLP_KV_REG_PCR_ENTRY_4_0                                                                    (32'h10018300)
`define KV_REG_PCR_ENTRY_4_0                                                                        (32'h300)
`define CLP_KV_REG_PCR_ENTRY_4_1                                                                    (32'h10018304)
`define KV_REG_PCR_ENTRY_4_1                                                                        (32'h304)
`define CLP_KV_REG_PCR_ENTRY_4_2                                                                    (32'h10018308)
`define KV_REG_PCR_ENTRY_4_2                                                                        (32'h308)
`define CLP_KV_REG_PCR_ENTRY_4_3                                                                    (32'h1001830c)
`define KV_REG_PCR_ENTRY_4_3                                                                        (32'h30c)
`define CLP_KV_REG_PCR_ENTRY_4_4                                                                    (32'h10018310)
`define KV_REG_PCR_ENTRY_4_4                                                                        (32'h310)
`define CLP_KV_REG_PCR_ENTRY_4_5                                                                    (32'h10018314)
`define KV_REG_PCR_ENTRY_4_5                                                                        (32'h314)
`define CLP_KV_REG_PCR_ENTRY_4_6                                                                    (32'h10018318)
`define KV_REG_PCR_ENTRY_4_6                                                                        (32'h318)
`define CLP_KV_REG_PCR_ENTRY_4_7                                                                    (32'h1001831c)
`define KV_REG_PCR_ENTRY_4_7                                                                        (32'h31c)
`define CLP_KV_REG_PCR_ENTRY_4_8                                                                    (32'h10018320)
`define KV_REG_PCR_ENTRY_4_8                                                                        (32'h320)
`define CLP_KV_REG_PCR_ENTRY_4_9                                                                    (32'h10018324)
`define KV_REG_PCR_ENTRY_4_9                                                                        (32'h324)
`define CLP_KV_REG_PCR_ENTRY_4_10                                                                   (32'h10018328)
`define KV_REG_PCR_ENTRY_4_10                                                                       (32'h328)
`define CLP_KV_REG_PCR_ENTRY_4_11                                                                   (32'h1001832c)
`define KV_REG_PCR_ENTRY_4_11                                                                       (32'h32c)
`define CLP_KV_REG_PCR_ENTRY_4_12                                                                   (32'h10018330)
`define KV_REG_PCR_ENTRY_4_12                                                                       (32'h330)
`define CLP_KV_REG_PCR_ENTRY_4_13                                                                   (32'h10018334)
`define KV_REG_PCR_ENTRY_4_13                                                                       (32'h334)
`define CLP_KV_REG_PCR_ENTRY_4_14                                                                   (32'h10018338)
`define KV_REG_PCR_ENTRY_4_14                                                                       (32'h338)
`define CLP_KV_REG_PCR_ENTRY_4_15                                                                   (32'h1001833c)
`define KV_REG_PCR_ENTRY_4_15                                                                       (32'h33c)
`define CLP_KV_REG_PCR_ENTRY_5_0                                                                    (32'h10018340)
`define KV_REG_PCR_ENTRY_5_0                                                                        (32'h340)
`define CLP_KV_REG_PCR_ENTRY_5_1                                                                    (32'h10018344)
`define KV_REG_PCR_ENTRY_5_1                                                                        (32'h344)
`define CLP_KV_REG_PCR_ENTRY_5_2                                                                    (32'h10018348)
`define KV_REG_PCR_ENTRY_5_2                                                                        (32'h348)
`define CLP_KV_REG_PCR_ENTRY_5_3                                                                    (32'h1001834c)
`define KV_REG_PCR_ENTRY_5_3                                                                        (32'h34c)
`define CLP_KV_REG_PCR_ENTRY_5_4                                                                    (32'h10018350)
`define KV_REG_PCR_ENTRY_5_4                                                                        (32'h350)
`define CLP_KV_REG_PCR_ENTRY_5_5                                                                    (32'h10018354)
`define KV_REG_PCR_ENTRY_5_5                                                                        (32'h354)
`define CLP_KV_REG_PCR_ENTRY_5_6                                                                    (32'h10018358)
`define KV_REG_PCR_ENTRY_5_6                                                                        (32'h358)
`define CLP_KV_REG_PCR_ENTRY_5_7                                                                    (32'h1001835c)
`define KV_REG_PCR_ENTRY_5_7                                                                        (32'h35c)
`define CLP_KV_REG_PCR_ENTRY_5_8                                                                    (32'h10018360)
`define KV_REG_PCR_ENTRY_5_8                                                                        (32'h360)
`define CLP_KV_REG_PCR_ENTRY_5_9                                                                    (32'h10018364)
`define KV_REG_PCR_ENTRY_5_9                                                                        (32'h364)
`define CLP_KV_REG_PCR_ENTRY_5_10                                                                   (32'h10018368)
`define KV_REG_PCR_ENTRY_5_10                                                                       (32'h368)
`define CLP_KV_REG_PCR_ENTRY_5_11                                                                   (32'h1001836c)
`define KV_REG_PCR_ENTRY_5_11                                                                       (32'h36c)
`define CLP_KV_REG_PCR_ENTRY_5_12                                                                   (32'h10018370)
`define KV_REG_PCR_ENTRY_5_12                                                                       (32'h370)
`define CLP_KV_REG_PCR_ENTRY_5_13                                                                   (32'h10018374)
`define KV_REG_PCR_ENTRY_5_13                                                                       (32'h374)
`define CLP_KV_REG_PCR_ENTRY_5_14                                                                   (32'h10018378)
`define KV_REG_PCR_ENTRY_5_14                                                                       (32'h378)
`define CLP_KV_REG_PCR_ENTRY_5_15                                                                   (32'h1001837c)
`define KV_REG_PCR_ENTRY_5_15                                                                       (32'h37c)
`define CLP_KV_REG_PCR_ENTRY_6_0                                                                    (32'h10018380)
`define KV_REG_PCR_ENTRY_6_0                                                                        (32'h380)
`define CLP_KV_REG_PCR_ENTRY_6_1                                                                    (32'h10018384)
`define KV_REG_PCR_ENTRY_6_1                                                                        (32'h384)
`define CLP_KV_REG_PCR_ENTRY_6_2                                                                    (32'h10018388)
`define KV_REG_PCR_ENTRY_6_2                                                                        (32'h388)
`define CLP_KV_REG_PCR_ENTRY_6_3                                                                    (32'h1001838c)
`define KV_REG_PCR_ENTRY_6_3                                                                        (32'h38c)
`define CLP_KV_REG_PCR_ENTRY_6_4                                                                    (32'h10018390)
`define KV_REG_PCR_ENTRY_6_4                                                                        (32'h390)
`define CLP_KV_REG_PCR_ENTRY_6_5                                                                    (32'h10018394)
`define KV_REG_PCR_ENTRY_6_5                                                                        (32'h394)
`define CLP_KV_REG_PCR_ENTRY_6_6                                                                    (32'h10018398)
`define KV_REG_PCR_ENTRY_6_6                                                                        (32'h398)
`define CLP_KV_REG_PCR_ENTRY_6_7                                                                    (32'h1001839c)
`define KV_REG_PCR_ENTRY_6_7                                                                        (32'h39c)
`define CLP_KV_REG_PCR_ENTRY_6_8                                                                    (32'h100183a0)
`define KV_REG_PCR_ENTRY_6_8                                                                        (32'h3a0)
`define CLP_KV_REG_PCR_ENTRY_6_9                                                                    (32'h100183a4)
`define KV_REG_PCR_ENTRY_6_9                                                                        (32'h3a4)
`define CLP_KV_REG_PCR_ENTRY_6_10                                                                   (32'h100183a8)
`define KV_REG_PCR_ENTRY_6_10                                                                       (32'h3a8)
`define CLP_KV_REG_PCR_ENTRY_6_11                                                                   (32'h100183ac)
`define KV_REG_PCR_ENTRY_6_11                                                                       (32'h3ac)
`define CLP_KV_REG_PCR_ENTRY_6_12                                                                   (32'h100183b0)
`define KV_REG_PCR_ENTRY_6_12                                                                       (32'h3b0)
`define CLP_KV_REG_PCR_ENTRY_6_13                                                                   (32'h100183b4)
`define KV_REG_PCR_ENTRY_6_13                                                                       (32'h3b4)
`define CLP_KV_REG_PCR_ENTRY_6_14                                                                   (32'h100183b8)
`define KV_REG_PCR_ENTRY_6_14                                                                       (32'h3b8)
`define CLP_KV_REG_PCR_ENTRY_6_15                                                                   (32'h100183bc)
`define KV_REG_PCR_ENTRY_6_15                                                                       (32'h3bc)
`define CLP_KV_REG_PCR_ENTRY_7_0                                                                    (32'h100183c0)
`define KV_REG_PCR_ENTRY_7_0                                                                        (32'h3c0)
`define CLP_KV_REG_PCR_ENTRY_7_1                                                                    (32'h100183c4)
`define KV_REG_PCR_ENTRY_7_1                                                                        (32'h3c4)
`define CLP_KV_REG_PCR_ENTRY_7_2                                                                    (32'h100183c8)
`define KV_REG_PCR_ENTRY_7_2                                                                        (32'h3c8)
`define CLP_KV_REG_PCR_ENTRY_7_3                                                                    (32'h100183cc)
`define KV_REG_PCR_ENTRY_7_3                                                                        (32'h3cc)
`define CLP_KV_REG_PCR_ENTRY_7_4                                                                    (32'h100183d0)
`define KV_REG_PCR_ENTRY_7_4                                                                        (32'h3d0)
`define CLP_KV_REG_PCR_ENTRY_7_5                                                                    (32'h100183d4)
`define KV_REG_PCR_ENTRY_7_5                                                                        (32'h3d4)
`define CLP_KV_REG_PCR_ENTRY_7_6                                                                    (32'h100183d8)
`define KV_REG_PCR_ENTRY_7_6                                                                        (32'h3d8)
`define CLP_KV_REG_PCR_ENTRY_7_7                                                                    (32'h100183dc)
`define KV_REG_PCR_ENTRY_7_7                                                                        (32'h3dc)
`define CLP_KV_REG_PCR_ENTRY_7_8                                                                    (32'h100183e0)
`define KV_REG_PCR_ENTRY_7_8                                                                        (32'h3e0)
`define CLP_KV_REG_PCR_ENTRY_7_9                                                                    (32'h100183e4)
`define KV_REG_PCR_ENTRY_7_9                                                                        (32'h3e4)
`define CLP_KV_REG_PCR_ENTRY_7_10                                                                   (32'h100183e8)
`define KV_REG_PCR_ENTRY_7_10                                                                       (32'h3e8)
`define CLP_KV_REG_PCR_ENTRY_7_11                                                                   (32'h100183ec)
`define KV_REG_PCR_ENTRY_7_11                                                                       (32'h3ec)
`define CLP_KV_REG_PCR_ENTRY_7_12                                                                   (32'h100183f0)
`define KV_REG_PCR_ENTRY_7_12                                                                       (32'h3f0)
`define CLP_KV_REG_PCR_ENTRY_7_13                                                                   (32'h100183f4)
`define KV_REG_PCR_ENTRY_7_13                                                                       (32'h3f4)
`define CLP_KV_REG_PCR_ENTRY_7_14                                                                   (32'h100183f8)
`define KV_REG_PCR_ENTRY_7_14                                                                       (32'h3f8)
`define CLP_KV_REG_PCR_ENTRY_7_15                                                                   (32'h100183fc)
`define KV_REG_PCR_ENTRY_7_15                                                                       (32'h3fc)
`define CLP_KV_REG_KEY_CTRL_0                                                                       (32'h10018400)
`define KV_REG_KEY_CTRL_0                                                                           (32'h400)
`define KV_REG_KEY_CTRL_0_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_0_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_0_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_0_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_0_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_0_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_0_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_0_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_0_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_0_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_KEY_CTRL_0_DEST_VALID_LOW                                                            (8)
`define KV_REG_KEY_CTRL_0_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_KEY_CTRL_0_RSVD_LOW                                                                  (14)
`define KV_REG_KEY_CTRL_0_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_KEY_CTRL_1                                                                       (32'h10018404)
`define KV_REG_KEY_CTRL_1                                                                           (32'h404)
`define KV_REG_KEY_CTRL_1_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_1_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_1_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_1_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_1_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_1_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_1_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_1_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_1_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_1_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_KEY_CTRL_1_DEST_VALID_LOW                                                            (8)
`define KV_REG_KEY_CTRL_1_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_KEY_CTRL_1_RSVD_LOW                                                                  (14)
`define KV_REG_KEY_CTRL_1_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_KEY_CTRL_2                                                                       (32'h10018408)
`define KV_REG_KEY_CTRL_2                                                                           (32'h408)
`define KV_REG_KEY_CTRL_2_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_2_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_2_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_2_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_2_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_2_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_2_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_2_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_2_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_2_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_KEY_CTRL_2_DEST_VALID_LOW                                                            (8)
`define KV_REG_KEY_CTRL_2_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_KEY_CTRL_2_RSVD_LOW                                                                  (14)
`define KV_REG_KEY_CTRL_2_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_KEY_CTRL_3                                                                       (32'h1001840c)
`define KV_REG_KEY_CTRL_3                                                                           (32'h40c)
`define KV_REG_KEY_CTRL_3_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_3_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_3_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_3_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_3_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_3_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_3_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_3_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_3_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_3_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_KEY_CTRL_3_DEST_VALID_LOW                                                            (8)
`define KV_REG_KEY_CTRL_3_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_KEY_CTRL_3_RSVD_LOW                                                                  (14)
`define KV_REG_KEY_CTRL_3_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_KEY_CTRL_4                                                                       (32'h10018410)
`define KV_REG_KEY_CTRL_4                                                                           (32'h410)
`define KV_REG_KEY_CTRL_4_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_4_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_4_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_4_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_4_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_4_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_4_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_4_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_4_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_4_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_KEY_CTRL_4_DEST_VALID_LOW                                                            (8)
`define KV_REG_KEY_CTRL_4_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_KEY_CTRL_4_RSVD_LOW                                                                  (14)
`define KV_REG_KEY_CTRL_4_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_KEY_CTRL_5                                                                       (32'h10018414)
`define KV_REG_KEY_CTRL_5                                                                           (32'h414)
`define KV_REG_KEY_CTRL_5_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_5_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_5_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_5_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_5_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_5_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_5_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_5_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_5_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_5_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_KEY_CTRL_5_DEST_VALID_LOW                                                            (8)
`define KV_REG_KEY_CTRL_5_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_KEY_CTRL_5_RSVD_LOW                                                                  (14)
`define KV_REG_KEY_CTRL_5_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_KEY_CTRL_6                                                                       (32'h10018418)
`define KV_REG_KEY_CTRL_6                                                                           (32'h418)
`define KV_REG_KEY_CTRL_6_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_6_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_6_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_6_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_6_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_6_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_6_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_6_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_6_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_6_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_KEY_CTRL_6_DEST_VALID_LOW                                                            (8)
`define KV_REG_KEY_CTRL_6_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_KEY_CTRL_6_RSVD_LOW                                                                  (14)
`define KV_REG_KEY_CTRL_6_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_KEY_CTRL_7                                                                       (32'h1001841c)
`define KV_REG_KEY_CTRL_7                                                                           (32'h41c)
`define KV_REG_KEY_CTRL_7_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_7_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_7_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_7_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_7_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_7_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_7_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_7_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_7_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_7_RSVD1_MASK                                                                (32'hf0)
`define KV_REG_KEY_CTRL_7_DEST_VALID_LOW                                                            (8)
`define KV_REG_KEY_CTRL_7_DEST_VALID_MASK                                                           (32'h3f00)
`define KV_REG_KEY_CTRL_7_RSVD_LOW                                                                  (14)
`define KV_REG_KEY_CTRL_7_RSVD_MASK                                                                 (32'hffffc000)
`define CLP_KV_REG_KEY_ENTRY_0_0                                                                    (32'h10018600)
`define KV_REG_KEY_ENTRY_0_0                                                                        (32'h600)
`define CLP_KV_REG_KEY_ENTRY_0_1                                                                    (32'h10018604)
`define KV_REG_KEY_ENTRY_0_1                                                                        (32'h604)
`define CLP_KV_REG_KEY_ENTRY_0_2                                                                    (32'h10018608)
`define KV_REG_KEY_ENTRY_0_2                                                                        (32'h608)
`define CLP_KV_REG_KEY_ENTRY_0_3                                                                    (32'h1001860c)
`define KV_REG_KEY_ENTRY_0_3                                                                        (32'h60c)
`define CLP_KV_REG_KEY_ENTRY_0_4                                                                    (32'h10018610)
`define KV_REG_KEY_ENTRY_0_4                                                                        (32'h610)
`define CLP_KV_REG_KEY_ENTRY_0_5                                                                    (32'h10018614)
`define KV_REG_KEY_ENTRY_0_5                                                                        (32'h614)
`define CLP_KV_REG_KEY_ENTRY_0_6                                                                    (32'h10018618)
`define KV_REG_KEY_ENTRY_0_6                                                                        (32'h618)
`define CLP_KV_REG_KEY_ENTRY_0_7                                                                    (32'h1001861c)
`define KV_REG_KEY_ENTRY_0_7                                                                        (32'h61c)
`define CLP_KV_REG_KEY_ENTRY_0_8                                                                    (32'h10018620)
`define KV_REG_KEY_ENTRY_0_8                                                                        (32'h620)
`define CLP_KV_REG_KEY_ENTRY_0_9                                                                    (32'h10018624)
`define KV_REG_KEY_ENTRY_0_9                                                                        (32'h624)
`define CLP_KV_REG_KEY_ENTRY_0_10                                                                   (32'h10018628)
`define KV_REG_KEY_ENTRY_0_10                                                                       (32'h628)
`define CLP_KV_REG_KEY_ENTRY_0_11                                                                   (32'h1001862c)
`define KV_REG_KEY_ENTRY_0_11                                                                       (32'h62c)
`define CLP_KV_REG_KEY_ENTRY_0_12                                                                   (32'h10018630)
`define KV_REG_KEY_ENTRY_0_12                                                                       (32'h630)
`define CLP_KV_REG_KEY_ENTRY_0_13                                                                   (32'h10018634)
`define KV_REG_KEY_ENTRY_0_13                                                                       (32'h634)
`define CLP_KV_REG_KEY_ENTRY_0_14                                                                   (32'h10018638)
`define KV_REG_KEY_ENTRY_0_14                                                                       (32'h638)
`define CLP_KV_REG_KEY_ENTRY_0_15                                                                   (32'h1001863c)
`define KV_REG_KEY_ENTRY_0_15                                                                       (32'h63c)
`define CLP_KV_REG_KEY_ENTRY_1_0                                                                    (32'h10018640)
`define KV_REG_KEY_ENTRY_1_0                                                                        (32'h640)
`define CLP_KV_REG_KEY_ENTRY_1_1                                                                    (32'h10018644)
`define KV_REG_KEY_ENTRY_1_1                                                                        (32'h644)
`define CLP_KV_REG_KEY_ENTRY_1_2                                                                    (32'h10018648)
`define KV_REG_KEY_ENTRY_1_2                                                                        (32'h648)
`define CLP_KV_REG_KEY_ENTRY_1_3                                                                    (32'h1001864c)
`define KV_REG_KEY_ENTRY_1_3                                                                        (32'h64c)
`define CLP_KV_REG_KEY_ENTRY_1_4                                                                    (32'h10018650)
`define KV_REG_KEY_ENTRY_1_4                                                                        (32'h650)
`define CLP_KV_REG_KEY_ENTRY_1_5                                                                    (32'h10018654)
`define KV_REG_KEY_ENTRY_1_5                                                                        (32'h654)
`define CLP_KV_REG_KEY_ENTRY_1_6                                                                    (32'h10018658)
`define KV_REG_KEY_ENTRY_1_6                                                                        (32'h658)
`define CLP_KV_REG_KEY_ENTRY_1_7                                                                    (32'h1001865c)
`define KV_REG_KEY_ENTRY_1_7                                                                        (32'h65c)
`define CLP_KV_REG_KEY_ENTRY_1_8                                                                    (32'h10018660)
`define KV_REG_KEY_ENTRY_1_8                                                                        (32'h660)
`define CLP_KV_REG_KEY_ENTRY_1_9                                                                    (32'h10018664)
`define KV_REG_KEY_ENTRY_1_9                                                                        (32'h664)
`define CLP_KV_REG_KEY_ENTRY_1_10                                                                   (32'h10018668)
`define KV_REG_KEY_ENTRY_1_10                                                                       (32'h668)
`define CLP_KV_REG_KEY_ENTRY_1_11                                                                   (32'h1001866c)
`define KV_REG_KEY_ENTRY_1_11                                                                       (32'h66c)
`define CLP_KV_REG_KEY_ENTRY_1_12                                                                   (32'h10018670)
`define KV_REG_KEY_ENTRY_1_12                                                                       (32'h670)
`define CLP_KV_REG_KEY_ENTRY_1_13                                                                   (32'h10018674)
`define KV_REG_KEY_ENTRY_1_13                                                                       (32'h674)
`define CLP_KV_REG_KEY_ENTRY_1_14                                                                   (32'h10018678)
`define KV_REG_KEY_ENTRY_1_14                                                                       (32'h678)
`define CLP_KV_REG_KEY_ENTRY_1_15                                                                   (32'h1001867c)
`define KV_REG_KEY_ENTRY_1_15                                                                       (32'h67c)
`define CLP_KV_REG_KEY_ENTRY_2_0                                                                    (32'h10018680)
`define KV_REG_KEY_ENTRY_2_0                                                                        (32'h680)
`define CLP_KV_REG_KEY_ENTRY_2_1                                                                    (32'h10018684)
`define KV_REG_KEY_ENTRY_2_1                                                                        (32'h684)
`define CLP_KV_REG_KEY_ENTRY_2_2                                                                    (32'h10018688)
`define KV_REG_KEY_ENTRY_2_2                                                                        (32'h688)
`define CLP_KV_REG_KEY_ENTRY_2_3                                                                    (32'h1001868c)
`define KV_REG_KEY_ENTRY_2_3                                                                        (32'h68c)
`define CLP_KV_REG_KEY_ENTRY_2_4                                                                    (32'h10018690)
`define KV_REG_KEY_ENTRY_2_4                                                                        (32'h690)
`define CLP_KV_REG_KEY_ENTRY_2_5                                                                    (32'h10018694)
`define KV_REG_KEY_ENTRY_2_5                                                                        (32'h694)
`define CLP_KV_REG_KEY_ENTRY_2_6                                                                    (32'h10018698)
`define KV_REG_KEY_ENTRY_2_6                                                                        (32'h698)
`define CLP_KV_REG_KEY_ENTRY_2_7                                                                    (32'h1001869c)
`define KV_REG_KEY_ENTRY_2_7                                                                        (32'h69c)
`define CLP_KV_REG_KEY_ENTRY_2_8                                                                    (32'h100186a0)
`define KV_REG_KEY_ENTRY_2_8                                                                        (32'h6a0)
`define CLP_KV_REG_KEY_ENTRY_2_9                                                                    (32'h100186a4)
`define KV_REG_KEY_ENTRY_2_9                                                                        (32'h6a4)
`define CLP_KV_REG_KEY_ENTRY_2_10                                                                   (32'h100186a8)
`define KV_REG_KEY_ENTRY_2_10                                                                       (32'h6a8)
`define CLP_KV_REG_KEY_ENTRY_2_11                                                                   (32'h100186ac)
`define KV_REG_KEY_ENTRY_2_11                                                                       (32'h6ac)
`define CLP_KV_REG_KEY_ENTRY_2_12                                                                   (32'h100186b0)
`define KV_REG_KEY_ENTRY_2_12                                                                       (32'h6b0)
`define CLP_KV_REG_KEY_ENTRY_2_13                                                                   (32'h100186b4)
`define KV_REG_KEY_ENTRY_2_13                                                                       (32'h6b4)
`define CLP_KV_REG_KEY_ENTRY_2_14                                                                   (32'h100186b8)
`define KV_REG_KEY_ENTRY_2_14                                                                       (32'h6b8)
`define CLP_KV_REG_KEY_ENTRY_2_15                                                                   (32'h100186bc)
`define KV_REG_KEY_ENTRY_2_15                                                                       (32'h6bc)
`define CLP_KV_REG_KEY_ENTRY_3_0                                                                    (32'h100186c0)
`define KV_REG_KEY_ENTRY_3_0                                                                        (32'h6c0)
`define CLP_KV_REG_KEY_ENTRY_3_1                                                                    (32'h100186c4)
`define KV_REG_KEY_ENTRY_3_1                                                                        (32'h6c4)
`define CLP_KV_REG_KEY_ENTRY_3_2                                                                    (32'h100186c8)
`define KV_REG_KEY_ENTRY_3_2                                                                        (32'h6c8)
`define CLP_KV_REG_KEY_ENTRY_3_3                                                                    (32'h100186cc)
`define KV_REG_KEY_ENTRY_3_3                                                                        (32'h6cc)
`define CLP_KV_REG_KEY_ENTRY_3_4                                                                    (32'h100186d0)
`define KV_REG_KEY_ENTRY_3_4                                                                        (32'h6d0)
`define CLP_KV_REG_KEY_ENTRY_3_5                                                                    (32'h100186d4)
`define KV_REG_KEY_ENTRY_3_5                                                                        (32'h6d4)
`define CLP_KV_REG_KEY_ENTRY_3_6                                                                    (32'h100186d8)
`define KV_REG_KEY_ENTRY_3_6                                                                        (32'h6d8)
`define CLP_KV_REG_KEY_ENTRY_3_7                                                                    (32'h100186dc)
`define KV_REG_KEY_ENTRY_3_7                                                                        (32'h6dc)
`define CLP_KV_REG_KEY_ENTRY_3_8                                                                    (32'h100186e0)
`define KV_REG_KEY_ENTRY_3_8                                                                        (32'h6e0)
`define CLP_KV_REG_KEY_ENTRY_3_9                                                                    (32'h100186e4)
`define KV_REG_KEY_ENTRY_3_9                                                                        (32'h6e4)
`define CLP_KV_REG_KEY_ENTRY_3_10                                                                   (32'h100186e8)
`define KV_REG_KEY_ENTRY_3_10                                                                       (32'h6e8)
`define CLP_KV_REG_KEY_ENTRY_3_11                                                                   (32'h100186ec)
`define KV_REG_KEY_ENTRY_3_11                                                                       (32'h6ec)
`define CLP_KV_REG_KEY_ENTRY_3_12                                                                   (32'h100186f0)
`define KV_REG_KEY_ENTRY_3_12                                                                       (32'h6f0)
`define CLP_KV_REG_KEY_ENTRY_3_13                                                                   (32'h100186f4)
`define KV_REG_KEY_ENTRY_3_13                                                                       (32'h6f4)
`define CLP_KV_REG_KEY_ENTRY_3_14                                                                   (32'h100186f8)
`define KV_REG_KEY_ENTRY_3_14                                                                       (32'h6f8)
`define CLP_KV_REG_KEY_ENTRY_3_15                                                                   (32'h100186fc)
`define KV_REG_KEY_ENTRY_3_15                                                                       (32'h6fc)
`define CLP_KV_REG_KEY_ENTRY_4_0                                                                    (32'h10018700)
`define KV_REG_KEY_ENTRY_4_0                                                                        (32'h700)
`define CLP_KV_REG_KEY_ENTRY_4_1                                                                    (32'h10018704)
`define KV_REG_KEY_ENTRY_4_1                                                                        (32'h704)
`define CLP_KV_REG_KEY_ENTRY_4_2                                                                    (32'h10018708)
`define KV_REG_KEY_ENTRY_4_2                                                                        (32'h708)
`define CLP_KV_REG_KEY_ENTRY_4_3                                                                    (32'h1001870c)
`define KV_REG_KEY_ENTRY_4_3                                                                        (32'h70c)
`define CLP_KV_REG_KEY_ENTRY_4_4                                                                    (32'h10018710)
`define KV_REG_KEY_ENTRY_4_4                                                                        (32'h710)
`define CLP_KV_REG_KEY_ENTRY_4_5                                                                    (32'h10018714)
`define KV_REG_KEY_ENTRY_4_5                                                                        (32'h714)
`define CLP_KV_REG_KEY_ENTRY_4_6                                                                    (32'h10018718)
`define KV_REG_KEY_ENTRY_4_6                                                                        (32'h718)
`define CLP_KV_REG_KEY_ENTRY_4_7                                                                    (32'h1001871c)
`define KV_REG_KEY_ENTRY_4_7                                                                        (32'h71c)
`define CLP_KV_REG_KEY_ENTRY_4_8                                                                    (32'h10018720)
`define KV_REG_KEY_ENTRY_4_8                                                                        (32'h720)
`define CLP_KV_REG_KEY_ENTRY_4_9                                                                    (32'h10018724)
`define KV_REG_KEY_ENTRY_4_9                                                                        (32'h724)
`define CLP_KV_REG_KEY_ENTRY_4_10                                                                   (32'h10018728)
`define KV_REG_KEY_ENTRY_4_10                                                                       (32'h728)
`define CLP_KV_REG_KEY_ENTRY_4_11                                                                   (32'h1001872c)
`define KV_REG_KEY_ENTRY_4_11                                                                       (32'h72c)
`define CLP_KV_REG_KEY_ENTRY_4_12                                                                   (32'h10018730)
`define KV_REG_KEY_ENTRY_4_12                                                                       (32'h730)
`define CLP_KV_REG_KEY_ENTRY_4_13                                                                   (32'h10018734)
`define KV_REG_KEY_ENTRY_4_13                                                                       (32'h734)
`define CLP_KV_REG_KEY_ENTRY_4_14                                                                   (32'h10018738)
`define KV_REG_KEY_ENTRY_4_14                                                                       (32'h738)
`define CLP_KV_REG_KEY_ENTRY_4_15                                                                   (32'h1001873c)
`define KV_REG_KEY_ENTRY_4_15                                                                       (32'h73c)
`define CLP_KV_REG_KEY_ENTRY_5_0                                                                    (32'h10018740)
`define KV_REG_KEY_ENTRY_5_0                                                                        (32'h740)
`define CLP_KV_REG_KEY_ENTRY_5_1                                                                    (32'h10018744)
`define KV_REG_KEY_ENTRY_5_1                                                                        (32'h744)
`define CLP_KV_REG_KEY_ENTRY_5_2                                                                    (32'h10018748)
`define KV_REG_KEY_ENTRY_5_2                                                                        (32'h748)
`define CLP_KV_REG_KEY_ENTRY_5_3                                                                    (32'h1001874c)
`define KV_REG_KEY_ENTRY_5_3                                                                        (32'h74c)
`define CLP_KV_REG_KEY_ENTRY_5_4                                                                    (32'h10018750)
`define KV_REG_KEY_ENTRY_5_4                                                                        (32'h750)
`define CLP_KV_REG_KEY_ENTRY_5_5                                                                    (32'h10018754)
`define KV_REG_KEY_ENTRY_5_5                                                                        (32'h754)
`define CLP_KV_REG_KEY_ENTRY_5_6                                                                    (32'h10018758)
`define KV_REG_KEY_ENTRY_5_6                                                                        (32'h758)
`define CLP_KV_REG_KEY_ENTRY_5_7                                                                    (32'h1001875c)
`define KV_REG_KEY_ENTRY_5_7                                                                        (32'h75c)
`define CLP_KV_REG_KEY_ENTRY_5_8                                                                    (32'h10018760)
`define KV_REG_KEY_ENTRY_5_8                                                                        (32'h760)
`define CLP_KV_REG_KEY_ENTRY_5_9                                                                    (32'h10018764)
`define KV_REG_KEY_ENTRY_5_9                                                                        (32'h764)
`define CLP_KV_REG_KEY_ENTRY_5_10                                                                   (32'h10018768)
`define KV_REG_KEY_ENTRY_5_10                                                                       (32'h768)
`define CLP_KV_REG_KEY_ENTRY_5_11                                                                   (32'h1001876c)
`define KV_REG_KEY_ENTRY_5_11                                                                       (32'h76c)
`define CLP_KV_REG_KEY_ENTRY_5_12                                                                   (32'h10018770)
`define KV_REG_KEY_ENTRY_5_12                                                                       (32'h770)
`define CLP_KV_REG_KEY_ENTRY_5_13                                                                   (32'h10018774)
`define KV_REG_KEY_ENTRY_5_13                                                                       (32'h774)
`define CLP_KV_REG_KEY_ENTRY_5_14                                                                   (32'h10018778)
`define KV_REG_KEY_ENTRY_5_14                                                                       (32'h778)
`define CLP_KV_REG_KEY_ENTRY_5_15                                                                   (32'h1001877c)
`define KV_REG_KEY_ENTRY_5_15                                                                       (32'h77c)
`define CLP_KV_REG_KEY_ENTRY_6_0                                                                    (32'h10018780)
`define KV_REG_KEY_ENTRY_6_0                                                                        (32'h780)
`define CLP_KV_REG_KEY_ENTRY_6_1                                                                    (32'h10018784)
`define KV_REG_KEY_ENTRY_6_1                                                                        (32'h784)
`define CLP_KV_REG_KEY_ENTRY_6_2                                                                    (32'h10018788)
`define KV_REG_KEY_ENTRY_6_2                                                                        (32'h788)
`define CLP_KV_REG_KEY_ENTRY_6_3                                                                    (32'h1001878c)
`define KV_REG_KEY_ENTRY_6_3                                                                        (32'h78c)
`define CLP_KV_REG_KEY_ENTRY_6_4                                                                    (32'h10018790)
`define KV_REG_KEY_ENTRY_6_4                                                                        (32'h790)
`define CLP_KV_REG_KEY_ENTRY_6_5                                                                    (32'h10018794)
`define KV_REG_KEY_ENTRY_6_5                                                                        (32'h794)
`define CLP_KV_REG_KEY_ENTRY_6_6                                                                    (32'h10018798)
`define KV_REG_KEY_ENTRY_6_6                                                                        (32'h798)
`define CLP_KV_REG_KEY_ENTRY_6_7                                                                    (32'h1001879c)
`define KV_REG_KEY_ENTRY_6_7                                                                        (32'h79c)
`define CLP_KV_REG_KEY_ENTRY_6_8                                                                    (32'h100187a0)
`define KV_REG_KEY_ENTRY_6_8                                                                        (32'h7a0)
`define CLP_KV_REG_KEY_ENTRY_6_9                                                                    (32'h100187a4)
`define KV_REG_KEY_ENTRY_6_9                                                                        (32'h7a4)
`define CLP_KV_REG_KEY_ENTRY_6_10                                                                   (32'h100187a8)
`define KV_REG_KEY_ENTRY_6_10                                                                       (32'h7a8)
`define CLP_KV_REG_KEY_ENTRY_6_11                                                                   (32'h100187ac)
`define KV_REG_KEY_ENTRY_6_11                                                                       (32'h7ac)
`define CLP_KV_REG_KEY_ENTRY_6_12                                                                   (32'h100187b0)
`define KV_REG_KEY_ENTRY_6_12                                                                       (32'h7b0)
`define CLP_KV_REG_KEY_ENTRY_6_13                                                                   (32'h100187b4)
`define KV_REG_KEY_ENTRY_6_13                                                                       (32'h7b4)
`define CLP_KV_REG_KEY_ENTRY_6_14                                                                   (32'h100187b8)
`define KV_REG_KEY_ENTRY_6_14                                                                       (32'h7b8)
`define CLP_KV_REG_KEY_ENTRY_6_15                                                                   (32'h100187bc)
`define KV_REG_KEY_ENTRY_6_15                                                                       (32'h7bc)
`define CLP_KV_REG_KEY_ENTRY_7_0                                                                    (32'h100187c0)
`define KV_REG_KEY_ENTRY_7_0                                                                        (32'h7c0)
`define CLP_KV_REG_KEY_ENTRY_7_1                                                                    (32'h100187c4)
`define KV_REG_KEY_ENTRY_7_1                                                                        (32'h7c4)
`define CLP_KV_REG_KEY_ENTRY_7_2                                                                    (32'h100187c8)
`define KV_REG_KEY_ENTRY_7_2                                                                        (32'h7c8)
`define CLP_KV_REG_KEY_ENTRY_7_3                                                                    (32'h100187cc)
`define KV_REG_KEY_ENTRY_7_3                                                                        (32'h7cc)
`define CLP_KV_REG_KEY_ENTRY_7_4                                                                    (32'h100187d0)
`define KV_REG_KEY_ENTRY_7_4                                                                        (32'h7d0)
`define CLP_KV_REG_KEY_ENTRY_7_5                                                                    (32'h100187d4)
`define KV_REG_KEY_ENTRY_7_5                                                                        (32'h7d4)
`define CLP_KV_REG_KEY_ENTRY_7_6                                                                    (32'h100187d8)
`define KV_REG_KEY_ENTRY_7_6                                                                        (32'h7d8)
`define CLP_KV_REG_KEY_ENTRY_7_7                                                                    (32'h100187dc)
`define KV_REG_KEY_ENTRY_7_7                                                                        (32'h7dc)
`define CLP_KV_REG_KEY_ENTRY_7_8                                                                    (32'h100187e0)
`define KV_REG_KEY_ENTRY_7_8                                                                        (32'h7e0)
`define CLP_KV_REG_KEY_ENTRY_7_9                                                                    (32'h100187e4)
`define KV_REG_KEY_ENTRY_7_9                                                                        (32'h7e4)
`define CLP_KV_REG_KEY_ENTRY_7_10                                                                   (32'h100187e8)
`define KV_REG_KEY_ENTRY_7_10                                                                       (32'h7e8)
`define CLP_KV_REG_KEY_ENTRY_7_11                                                                   (32'h100187ec)
`define KV_REG_KEY_ENTRY_7_11                                                                       (32'h7ec)
`define CLP_KV_REG_KEY_ENTRY_7_12                                                                   (32'h100187f0)
`define KV_REG_KEY_ENTRY_7_12                                                                       (32'h7f0)
`define CLP_KV_REG_KEY_ENTRY_7_13                                                                   (32'h100187f4)
`define KV_REG_KEY_ENTRY_7_13                                                                       (32'h7f4)
`define CLP_KV_REG_KEY_ENTRY_7_14                                                                   (32'h100187f8)
`define KV_REG_KEY_ENTRY_7_14                                                                       (32'h7f8)
`define CLP_KV_REG_KEY_ENTRY_7_15                                                                   (32'h100187fc)
`define KV_REG_KEY_ENTRY_7_15                                                                       (32'h7fc)
`define CLP_KV_REG_CLEAR_SECRETS                                                                    (32'h10018800)
`define KV_REG_CLEAR_SECRETS                                                                        (32'h800)
`define KV_REG_CLEAR_SECRETS_WR_DEBUG_VALUES_LOW                                                    (0)
`define KV_REG_CLEAR_SECRETS_WR_DEBUG_VALUES_MASK                                                   (32'h1)
`define KV_REG_CLEAR_SECRETS_SEL_DEBUG_VALUE_LOW                                                    (1)
`define KV_REG_CLEAR_SECRETS_SEL_DEBUG_VALUE_MASK                                                   (32'h2)
`define CLP_SHA512_REG_BASE_ADDR                                                                    (32'h10020000)
`define CLP_SHA512_REG_SHA512_NAME_0                                                                (32'h10020000)
`define SHA512_REG_SHA512_NAME_0                                                                    (32'h0)
`define CLP_SHA512_REG_SHA512_NAME_1                                                                (32'h10020004)
`define SHA512_REG_SHA512_NAME_1                                                                    (32'h4)
`define CLP_SHA512_REG_SHA512_VERSION_0                                                             (32'h10020008)
`define SHA512_REG_SHA512_VERSION_0                                                                 (32'h8)
`define CLP_SHA512_REG_SHA512_VERSION_1                                                             (32'h1002000c)
`define SHA512_REG_SHA512_VERSION_1                                                                 (32'hc)
`define CLP_SHA512_REG_SHA512_CTRL                                                                  (32'h10020010)
`define SHA512_REG_SHA512_CTRL                                                                      (32'h10)
`define SHA512_REG_SHA512_CTRL_INIT_LOW                                                             (0)
`define SHA512_REG_SHA512_CTRL_INIT_MASK                                                            (32'h1)
`define SHA512_REG_SHA512_CTRL_NEXT_LOW                                                             (1)
`define SHA512_REG_SHA512_CTRL_NEXT_MASK                                                            (32'h2)
`define SHA512_REG_SHA512_CTRL_MODE_LOW                                                             (2)
`define SHA512_REG_SHA512_CTRL_MODE_MASK                                                            (32'hc)
`define SHA512_REG_SHA512_CTRL_ZEROIZE_LOW                                                          (4)
`define SHA512_REG_SHA512_CTRL_ZEROIZE_MASK                                                         (32'h10)
`define CLP_SHA512_REG_SHA512_STATUS                                                                (32'h10020018)
`define SHA512_REG_SHA512_STATUS                                                                    (32'h18)
`define SHA512_REG_SHA512_STATUS_READY_LOW                                                          (0)
`define SHA512_REG_SHA512_STATUS_READY_MASK                                                         (32'h1)
`define SHA512_REG_SHA512_STATUS_VALID_LOW                                                          (1)
`define SHA512_REG_SHA512_STATUS_VALID_MASK                                                         (32'h2)
`define CLP_SHA512_REG_SHA512_BLOCK_0                                                               (32'h10020080)
`define SHA512_REG_SHA512_BLOCK_0                                                                   (32'h80)
`define CLP_SHA512_REG_SHA512_BLOCK_1                                                               (32'h10020084)
`define SHA512_REG_SHA512_BLOCK_1                                                                   (32'h84)
`define CLP_SHA512_REG_SHA512_BLOCK_2                                                               (32'h10020088)
`define SHA512_REG_SHA512_BLOCK_2                                                                   (32'h88)
`define CLP_SHA512_REG_SHA512_BLOCK_3                                                               (32'h1002008c)
`define SHA512_REG_SHA512_BLOCK_3                                                                   (32'h8c)
`define CLP_SHA512_REG_SHA512_BLOCK_4                                                               (32'h10020090)
`define SHA512_REG_SHA512_BLOCK_4                                                                   (32'h90)
`define CLP_SHA512_REG_SHA512_BLOCK_5                                                               (32'h10020094)
`define SHA512_REG_SHA512_BLOCK_5                                                                   (32'h94)
`define CLP_SHA512_REG_SHA512_BLOCK_6                                                               (32'h10020098)
`define SHA512_REG_SHA512_BLOCK_6                                                                   (32'h98)
`define CLP_SHA512_REG_SHA512_BLOCK_7                                                               (32'h1002009c)
`define SHA512_REG_SHA512_BLOCK_7                                                                   (32'h9c)
`define CLP_SHA512_REG_SHA512_BLOCK_8                                                               (32'h100200a0)
`define SHA512_REG_SHA512_BLOCK_8                                                                   (32'ha0)
`define CLP_SHA512_REG_SHA512_BLOCK_9                                                               (32'h100200a4)
`define SHA512_REG_SHA512_BLOCK_9                                                                   (32'ha4)
`define CLP_SHA512_REG_SHA512_BLOCK_10                                                              (32'h100200a8)
`define SHA512_REG_SHA512_BLOCK_10                                                                  (32'ha8)
`define CLP_SHA512_REG_SHA512_BLOCK_11                                                              (32'h100200ac)
`define SHA512_REG_SHA512_BLOCK_11                                                                  (32'hac)
`define CLP_SHA512_REG_SHA512_BLOCK_12                                                              (32'h100200b0)
`define SHA512_REG_SHA512_BLOCK_12                                                                  (32'hb0)
`define CLP_SHA512_REG_SHA512_BLOCK_13                                                              (32'h100200b4)
`define SHA512_REG_SHA512_BLOCK_13                                                                  (32'hb4)
`define CLP_SHA512_REG_SHA512_BLOCK_14                                                              (32'h100200b8)
`define SHA512_REG_SHA512_BLOCK_14                                                                  (32'hb8)
`define CLP_SHA512_REG_SHA512_BLOCK_15                                                              (32'h100200bc)
`define SHA512_REG_SHA512_BLOCK_15                                                                  (32'hbc)
`define CLP_SHA512_REG_SHA512_BLOCK_16                                                              (32'h100200c0)
`define SHA512_REG_SHA512_BLOCK_16                                                                  (32'hc0)
`define CLP_SHA512_REG_SHA512_BLOCK_17                                                              (32'h100200c4)
`define SHA512_REG_SHA512_BLOCK_17                                                                  (32'hc4)
`define CLP_SHA512_REG_SHA512_BLOCK_18                                                              (32'h100200c8)
`define SHA512_REG_SHA512_BLOCK_18                                                                  (32'hc8)
`define CLP_SHA512_REG_SHA512_BLOCK_19                                                              (32'h100200cc)
`define SHA512_REG_SHA512_BLOCK_19                                                                  (32'hcc)
`define CLP_SHA512_REG_SHA512_BLOCK_20                                                              (32'h100200d0)
`define SHA512_REG_SHA512_BLOCK_20                                                                  (32'hd0)
`define CLP_SHA512_REG_SHA512_BLOCK_21                                                              (32'h100200d4)
`define SHA512_REG_SHA512_BLOCK_21                                                                  (32'hd4)
`define CLP_SHA512_REG_SHA512_BLOCK_22                                                              (32'h100200d8)
`define SHA512_REG_SHA512_BLOCK_22                                                                  (32'hd8)
`define CLP_SHA512_REG_SHA512_BLOCK_23                                                              (32'h100200dc)
`define SHA512_REG_SHA512_BLOCK_23                                                                  (32'hdc)
`define CLP_SHA512_REG_SHA512_BLOCK_24                                                              (32'h100200e0)
`define SHA512_REG_SHA512_BLOCK_24                                                                  (32'he0)
`define CLP_SHA512_REG_SHA512_BLOCK_25                                                              (32'h100200e4)
`define SHA512_REG_SHA512_BLOCK_25                                                                  (32'he4)
`define CLP_SHA512_REG_SHA512_BLOCK_26                                                              (32'h100200e8)
`define SHA512_REG_SHA512_BLOCK_26                                                                  (32'he8)
`define CLP_SHA512_REG_SHA512_BLOCK_27                                                              (32'h100200ec)
`define SHA512_REG_SHA512_BLOCK_27                                                                  (32'hec)
`define CLP_SHA512_REG_SHA512_BLOCK_28                                                              (32'h100200f0)
`define SHA512_REG_SHA512_BLOCK_28                                                                  (32'hf0)
`define CLP_SHA512_REG_SHA512_BLOCK_29                                                              (32'h100200f4)
`define SHA512_REG_SHA512_BLOCK_29                                                                  (32'hf4)
`define CLP_SHA512_REG_SHA512_BLOCK_30                                                              (32'h100200f8)
`define SHA512_REG_SHA512_BLOCK_30                                                                  (32'hf8)
`define CLP_SHA512_REG_SHA512_BLOCK_31                                                              (32'h100200fc)
`define SHA512_REG_SHA512_BLOCK_31                                                                  (32'hfc)
`define CLP_SHA512_REG_SHA512_DIGEST_0                                                              (32'h10020100)
`define SHA512_REG_SHA512_DIGEST_0                                                                  (32'h100)
`define CLP_SHA512_REG_SHA512_DIGEST_1                                                              (32'h10020104)
`define SHA512_REG_SHA512_DIGEST_1                                                                  (32'h104)
`define CLP_SHA512_REG_SHA512_DIGEST_2                                                              (32'h10020108)
`define SHA512_REG_SHA512_DIGEST_2                                                                  (32'h108)
`define CLP_SHA512_REG_SHA512_DIGEST_3                                                              (32'h1002010c)
`define SHA512_REG_SHA512_DIGEST_3                                                                  (32'h10c)
`define CLP_SHA512_REG_SHA512_DIGEST_4                                                              (32'h10020110)
`define SHA512_REG_SHA512_DIGEST_4                                                                  (32'h110)
`define CLP_SHA512_REG_SHA512_DIGEST_5                                                              (32'h10020114)
`define SHA512_REG_SHA512_DIGEST_5                                                                  (32'h114)
`define CLP_SHA512_REG_SHA512_DIGEST_6                                                              (32'h10020118)
`define SHA512_REG_SHA512_DIGEST_6                                                                  (32'h118)
`define CLP_SHA512_REG_SHA512_DIGEST_7                                                              (32'h1002011c)
`define SHA512_REG_SHA512_DIGEST_7                                                                  (32'h11c)
`define CLP_SHA512_REG_SHA512_DIGEST_8                                                              (32'h10020120)
`define SHA512_REG_SHA512_DIGEST_8                                                                  (32'h120)
`define CLP_SHA512_REG_SHA512_DIGEST_9                                                              (32'h10020124)
`define SHA512_REG_SHA512_DIGEST_9                                                                  (32'h124)
`define CLP_SHA512_REG_SHA512_DIGEST_10                                                             (32'h10020128)
`define SHA512_REG_SHA512_DIGEST_10                                                                 (32'h128)
`define CLP_SHA512_REG_SHA512_DIGEST_11                                                             (32'h1002012c)
`define SHA512_REG_SHA512_DIGEST_11                                                                 (32'h12c)
`define CLP_SHA512_REG_SHA512_DIGEST_12                                                             (32'h10020130)
`define SHA512_REG_SHA512_DIGEST_12                                                                 (32'h130)
`define CLP_SHA512_REG_SHA512_DIGEST_13                                                             (32'h10020134)
`define SHA512_REG_SHA512_DIGEST_13                                                                 (32'h134)
`define CLP_SHA512_REG_SHA512_DIGEST_14                                                             (32'h10020138)
`define SHA512_REG_SHA512_DIGEST_14                                                                 (32'h138)
`define CLP_SHA512_REG_SHA512_DIGEST_15                                                             (32'h1002013c)
`define SHA512_REG_SHA512_DIGEST_15                                                                 (32'h13c)
`define CLP_SHA512_REG_SHA512_KV_RD_CTRL                                                            (32'h10020600)
`define SHA512_REG_SHA512_KV_RD_CTRL                                                                (32'h600)
`define SHA512_REG_SHA512_KV_RD_CTRL_READ_EN_LOW                                                    (0)
`define SHA512_REG_SHA512_KV_RD_CTRL_READ_EN_MASK                                                   (32'h1)
`define SHA512_REG_SHA512_KV_RD_CTRL_READ_ENTRY_LOW                                                 (1)
`define SHA512_REG_SHA512_KV_RD_CTRL_READ_ENTRY_MASK                                                (32'he)
`define SHA512_REG_SHA512_KV_RD_CTRL_ENTRY_IS_PCR_LOW                                               (4)
`define SHA512_REG_SHA512_KV_RD_CTRL_ENTRY_IS_PCR_MASK                                              (32'h10)
`define SHA512_REG_SHA512_KV_RD_CTRL_ENTRY_DATA_SIZE_LOW                                            (5)
`define SHA512_REG_SHA512_KV_RD_CTRL_ENTRY_DATA_SIZE_MASK                                           (32'h3e0)
`define SHA512_REG_SHA512_KV_RD_CTRL_RSVD_LOW                                                       (10)
`define SHA512_REG_SHA512_KV_RD_CTRL_RSVD_MASK                                                      (32'h3ffffc00)
`define CLP_SHA512_REG_SHA512_KV_RD_STATUS                                                          (32'h10020604)
`define SHA512_REG_SHA512_KV_RD_STATUS                                                              (32'h604)
`define SHA512_REG_SHA512_KV_RD_STATUS_READY_LOW                                                    (0)
`define SHA512_REG_SHA512_KV_RD_STATUS_READY_MASK                                                   (32'h1)
`define SHA512_REG_SHA512_KV_RD_STATUS_VALID_LOW                                                    (1)
`define SHA512_REG_SHA512_KV_RD_STATUS_VALID_MASK                                                   (32'h2)
`define SHA512_REG_SHA512_KV_RD_STATUS_ERROR_LOW                                                    (2)
`define SHA512_REG_SHA512_KV_RD_STATUS_ERROR_MASK                                                   (32'h3fc)
`define CLP_SHA512_REG_SHA512_KV_WR_CTRL                                                            (32'h10020608)
`define SHA512_REG_SHA512_KV_WR_CTRL                                                                (32'h608)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_EN_LOW                                                   (0)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_EN_MASK                                                  (32'h1)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_ENTRY_LOW                                                (1)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_ENTRY_MASK                                               (32'he)
`define SHA512_REG_SHA512_KV_WR_CTRL_ENTRY_IS_PCR_LOW                                               (4)
`define SHA512_REG_SHA512_KV_WR_CTRL_ENTRY_IS_PCR_MASK                                              (32'h10)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_KEY_DEST_VALID_LOW                                        (5)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_KEY_DEST_VALID_MASK                                       (32'h20)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                      (6)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                     (32'h40)
`define SHA512_REG_SHA512_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_LOW                                       (7)
`define SHA512_REG_SHA512_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_MASK                                      (32'h80)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_PKEY_DEST_VALID_LOW                                        (8)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_PKEY_DEST_VALID_MASK                                       (32'h100)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_SEED_DEST_VALID_LOW                                        (9)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_SEED_DEST_VALID_MASK                                       (32'h200)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_MSG_DEST_VALID_LOW                                         (10)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_MSG_DEST_VALID_MASK                                        (32'h400)
`define SHA512_REG_SHA512_KV_WR_CTRL_RSVD_LOW                                                       (11)
`define SHA512_REG_SHA512_KV_WR_CTRL_RSVD_MASK                                                      (32'h3ffff800)
`define CLP_SHA512_REG_SHA512_KV_WR_STATUS                                                          (32'h1002060c)
`define SHA512_REG_SHA512_KV_WR_STATUS                                                              (32'h60c)
`define SHA512_REG_SHA512_KV_WR_STATUS_READY_LOW                                                    (0)
`define SHA512_REG_SHA512_KV_WR_STATUS_READY_MASK                                                   (32'h1)
`define SHA512_REG_SHA512_KV_WR_STATUS_VALID_LOW                                                    (1)
`define SHA512_REG_SHA512_KV_WR_STATUS_VALID_MASK                                                   (32'h2)
`define SHA512_REG_SHA512_KV_WR_STATUS_ERROR_LOW                                                    (2)
`define SHA512_REG_SHA512_KV_WR_STATUS_ERROR_MASK                                                   (32'h3fc)
`define CLP_SHA512_REG_INTR_BLOCK_RF_START                                                          (32'h10020800)
`define CLP_SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h10020800)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                   (32'h800)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                      (0)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                     (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                      (1)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                     (32'h2)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h10020804)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                    (32'h804)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                      (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                     (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                      (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                     (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                      (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                     (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                      (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                     (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h10020808)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                    (32'h808)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                              (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                             (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h1002080c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                (32'h80c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h10020810)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                (32'h810)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h10020814)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                              (32'h814)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                               (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                              (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                               (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                              (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                               (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                              (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                               (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                              (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h10020818)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                              (32'h818)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                       (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                      (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h1002081c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                  (32'h81c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                  (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                 (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                  (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                 (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                  (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                 (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                  (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                 (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h10020820)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                  (32'h820)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                          (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                         (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h10020900)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                (32'h900)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h10020904)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                (32'h904)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h10020908)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                (32'h908)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h1002090c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                (32'h90c)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h10020980)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                        (32'h980)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'h10020a00)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                           (32'ha00)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'h10020a04)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                           (32'ha04)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'h10020a08)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                           (32'ha08)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'h10020a0c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                           (32'ha0c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'h10020a10)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                   (32'ha10)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_SHA256_REG_BASE_ADDR                                                                    (32'h10028000)
`define CLP_SHA256_REG_SHA256_NAME_0                                                                (32'h10028000)
`define SHA256_REG_SHA256_NAME_0                                                                    (32'h0)
`define CLP_SHA256_REG_SHA256_NAME_1                                                                (32'h10028004)
`define SHA256_REG_SHA256_NAME_1                                                                    (32'h4)
`define CLP_SHA256_REG_SHA256_VERSION_0                                                             (32'h10028008)
`define SHA256_REG_SHA256_VERSION_0                                                                 (32'h8)
`define CLP_SHA256_REG_SHA256_VERSION_1                                                             (32'h1002800c)
`define SHA256_REG_SHA256_VERSION_1                                                                 (32'hc)
`define CLP_SHA256_REG_SHA256_CTRL                                                                  (32'h10028010)
`define SHA256_REG_SHA256_CTRL                                                                      (32'h10)
`define SHA256_REG_SHA256_CTRL_INIT_LOW                                                             (0)
`define SHA256_REG_SHA256_CTRL_INIT_MASK                                                            (32'h1)
`define SHA256_REG_SHA256_CTRL_NEXT_LOW                                                             (1)
`define SHA256_REG_SHA256_CTRL_NEXT_MASK                                                            (32'h2)
`define SHA256_REG_SHA256_CTRL_MODE_LOW                                                             (2)
`define SHA256_REG_SHA256_CTRL_MODE_MASK                                                            (32'h4)
`define CLP_SHA256_REG_SHA256_STATUS                                                                (32'h10028018)
`define SHA256_REG_SHA256_STATUS                                                                    (32'h18)
`define SHA256_REG_SHA256_STATUS_READY_LOW                                                          (0)
`define SHA256_REG_SHA256_STATUS_READY_MASK                                                         (32'h1)
`define SHA256_REG_SHA256_STATUS_VALID_LOW                                                          (1)
`define SHA256_REG_SHA256_STATUS_VALID_MASK                                                         (32'h2)
`define CLP_SHA256_REG_SHA256_BLOCK_0                                                               (32'h10028080)
`define SHA256_REG_SHA256_BLOCK_0                                                                   (32'h80)
`define CLP_SHA256_REG_SHA256_BLOCK_1                                                               (32'h10028084)
`define SHA256_REG_SHA256_BLOCK_1                                                                   (32'h84)
`define CLP_SHA256_REG_SHA256_BLOCK_2                                                               (32'h10028088)
`define SHA256_REG_SHA256_BLOCK_2                                                                   (32'h88)
`define CLP_SHA256_REG_SHA256_BLOCK_3                                                               (32'h1002808c)
`define SHA256_REG_SHA256_BLOCK_3                                                                   (32'h8c)
`define CLP_SHA256_REG_SHA256_BLOCK_4                                                               (32'h10028090)
`define SHA256_REG_SHA256_BLOCK_4                                                                   (32'h90)
`define CLP_SHA256_REG_SHA256_BLOCK_5                                                               (32'h10028094)
`define SHA256_REG_SHA256_BLOCK_5                                                                   (32'h94)
`define CLP_SHA256_REG_SHA256_BLOCK_6                                                               (32'h10028098)
`define SHA256_REG_SHA256_BLOCK_6                                                                   (32'h98)
`define CLP_SHA256_REG_SHA256_BLOCK_7                                                               (32'h1002809c)
`define SHA256_REG_SHA256_BLOCK_7                                                                   (32'h9c)
`define CLP_SHA256_REG_SHA256_BLOCK_8                                                               (32'h100280a0)
`define SHA256_REG_SHA256_BLOCK_8                                                                   (32'ha0)
`define CLP_SHA256_REG_SHA256_BLOCK_9                                                               (32'h100280a4)
`define SHA256_REG_SHA256_BLOCK_9                                                                   (32'ha4)
`define CLP_SHA256_REG_SHA256_BLOCK_10                                                              (32'h100280a8)
`define SHA256_REG_SHA256_BLOCK_10                                                                  (32'ha8)
`define CLP_SHA256_REG_SHA256_BLOCK_11                                                              (32'h100280ac)
`define SHA256_REG_SHA256_BLOCK_11                                                                  (32'hac)
`define CLP_SHA256_REG_SHA256_BLOCK_12                                                              (32'h100280b0)
`define SHA256_REG_SHA256_BLOCK_12                                                                  (32'hb0)
`define CLP_SHA256_REG_SHA256_BLOCK_13                                                              (32'h100280b4)
`define SHA256_REG_SHA256_BLOCK_13                                                                  (32'hb4)
`define CLP_SHA256_REG_SHA256_BLOCK_14                                                              (32'h100280b8)
`define SHA256_REG_SHA256_BLOCK_14                                                                  (32'hb8)
`define CLP_SHA256_REG_SHA256_BLOCK_15                                                              (32'h100280bc)
`define SHA256_REG_SHA256_BLOCK_15                                                                  (32'hbc)
`define CLP_SHA256_REG_SHA256_DIGEST_0                                                              (32'h10028100)
`define SHA256_REG_SHA256_DIGEST_0                                                                  (32'h100)
`define CLP_SHA256_REG_SHA256_DIGEST_1                                                              (32'h10028104)
`define SHA256_REG_SHA256_DIGEST_1                                                                  (32'h104)
`define CLP_SHA256_REG_SHA256_DIGEST_2                                                              (32'h10028108)
`define SHA256_REG_SHA256_DIGEST_2                                                                  (32'h108)
`define CLP_SHA256_REG_SHA256_DIGEST_3                                                              (32'h1002810c)
`define SHA256_REG_SHA256_DIGEST_3                                                                  (32'h10c)
`define CLP_SHA256_REG_SHA256_DIGEST_4                                                              (32'h10028110)
`define SHA256_REG_SHA256_DIGEST_4                                                                  (32'h110)
`define CLP_SHA256_REG_SHA256_DIGEST_5                                                              (32'h10028114)
`define SHA256_REG_SHA256_DIGEST_5                                                                  (32'h114)
`define CLP_SHA256_REG_SHA256_DIGEST_6                                                              (32'h10028118)
`define SHA256_REG_SHA256_DIGEST_6                                                                  (32'h118)
`define CLP_SHA256_REG_SHA256_DIGEST_7                                                              (32'h1002811c)
`define SHA256_REG_SHA256_DIGEST_7                                                                  (32'h11c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_START                                                          (32'h10028800)
`define CLP_SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h10028800)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                   (32'h800)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                      (0)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                     (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                      (1)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                     (32'h2)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h10028804)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                    (32'h804)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                      (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                     (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                      (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                     (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                      (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                     (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                      (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                     (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h10028808)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                    (32'h808)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                              (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                             (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h1002880c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                (32'h80c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h10028810)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                (32'h810)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h10028814)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                              (32'h814)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                               (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                              (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                               (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                              (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                               (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                              (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                               (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                              (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h10028818)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                              (32'h818)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                       (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                      (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h1002881c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                  (32'h81c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                  (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                 (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                  (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                 (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                  (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                 (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                  (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                 (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h10028820)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                  (32'h820)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                          (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                         (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h10028900)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                (32'h900)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h10028904)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                (32'h904)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h10028908)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                (32'h908)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h1002890c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                (32'h90c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h10028980)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                        (32'h980)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'h10028a00)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                           (32'ha00)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'h10028a04)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                           (32'ha04)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'h10028a08)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                           (32'ha08)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'h10028a0c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                           (32'ha0c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'h10028a10)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                   (32'ha10)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_MBOX_CSR_BASE_ADDR                                                                      (32'h30020000)
`define CLP_MBOX_CSR_MBOX_LOCK                                                                      (32'h30020000)
`define MBOX_CSR_MBOX_LOCK                                                                          (32'h0)
`define MBOX_CSR_MBOX_LOCK_LOCK_LOW                                                                 (0)
`define MBOX_CSR_MBOX_LOCK_LOCK_MASK                                                                (32'h1)
`define CLP_MBOX_CSR_MBOX_USER                                                                      (32'h30020004)
`define MBOX_CSR_MBOX_USER                                                                          (32'h4)
`define CLP_MBOX_CSR_MBOX_CMD                                                                       (32'h30020008)
`define MBOX_CSR_MBOX_CMD                                                                           (32'h8)
`define CLP_MBOX_CSR_MBOX_DLEN                                                                      (32'h3002000c)
`define MBOX_CSR_MBOX_DLEN                                                                          (32'hc)
`define CLP_MBOX_CSR_MBOX_DATAIN                                                                    (32'h30020010)
`define MBOX_CSR_MBOX_DATAIN                                                                        (32'h10)
`define CLP_MBOX_CSR_MBOX_DATAOUT                                                                   (32'h30020014)
`define MBOX_CSR_MBOX_DATAOUT                                                                       (32'h14)
`define CLP_MBOX_CSR_MBOX_EXECUTE                                                                   (32'h30020018)
`define MBOX_CSR_MBOX_EXECUTE                                                                       (32'h18)
`define MBOX_CSR_MBOX_EXECUTE_EXECUTE_LOW                                                           (0)
`define MBOX_CSR_MBOX_EXECUTE_EXECUTE_MASK                                                          (32'h1)
`define CLP_MBOX_CSR_MBOX_STATUS                                                                    (32'h3002001c)
`define MBOX_CSR_MBOX_STATUS                                                                        (32'h1c)
`define MBOX_CSR_MBOX_STATUS_STATUS_LOW                                                             (0)
`define MBOX_CSR_MBOX_STATUS_STATUS_MASK                                                            (32'hf)
`define MBOX_CSR_MBOX_STATUS_ECC_SINGLE_ERROR_LOW                                                   (4)
`define MBOX_CSR_MBOX_STATUS_ECC_SINGLE_ERROR_MASK                                                  (32'h10)
`define MBOX_CSR_MBOX_STATUS_ECC_DOUBLE_ERROR_LOW                                                   (5)
`define MBOX_CSR_MBOX_STATUS_ECC_DOUBLE_ERROR_MASK                                                  (32'h20)
`define MBOX_CSR_MBOX_STATUS_MBOX_FSM_PS_LOW                                                        (6)
`define MBOX_CSR_MBOX_STATUS_MBOX_FSM_PS_MASK                                                       (32'h1c0)
`define MBOX_CSR_MBOX_STATUS_SOC_HAS_LOCK_LOW                                                       (9)
`define MBOX_CSR_MBOX_STATUS_SOC_HAS_LOCK_MASK                                                      (32'h200)
`define CLP_MBOX_CSR_MBOX_UNLOCK                                                                    (32'h30020020)
`define MBOX_CSR_MBOX_UNLOCK                                                                        (32'h20)
`define MBOX_CSR_MBOX_UNLOCK_UNLOCK_LOW                                                             (0)
`define MBOX_CSR_MBOX_UNLOCK_UNLOCK_MASK                                                            (32'h1)
`define CLP_SHA512_ACC_CSR_BASE_ADDR                                                                (32'h30021000)
`define CLP_SHA512_ACC_CSR_LOCK                                                                     (32'h30021000)
`define SHA512_ACC_CSR_LOCK                                                                         (32'h0)
`define SHA512_ACC_CSR_LOCK_LOCK_LOW                                                                (0)
`define SHA512_ACC_CSR_LOCK_LOCK_MASK                                                               (32'h1)
`define CLP_SHA512_ACC_CSR_USER                                                                     (32'h30021004)
`define SHA512_ACC_CSR_USER                                                                         (32'h4)
`define CLP_SHA512_ACC_CSR_MODE                                                                     (32'h30021008)
`define SHA512_ACC_CSR_MODE                                                                         (32'h8)
`define SHA512_ACC_CSR_MODE_MODE_LOW                                                                (0)
`define SHA512_ACC_CSR_MODE_MODE_MASK                                                               (32'h3)
`define SHA512_ACC_CSR_MODE_ENDIAN_TOGGLE_LOW                                                       (2)
`define SHA512_ACC_CSR_MODE_ENDIAN_TOGGLE_MASK                                                      (32'h4)
`define CLP_SHA512_ACC_CSR_START_ADDRESS                                                            (32'h3002100c)
`define SHA512_ACC_CSR_START_ADDRESS                                                                (32'hc)
`define CLP_SHA512_ACC_CSR_DLEN                                                                     (32'h30021010)
`define SHA512_ACC_CSR_DLEN                                                                         (32'h10)
`define CLP_SHA512_ACC_CSR_DATAIN                                                                   (32'h30021014)
`define SHA512_ACC_CSR_DATAIN                                                                       (32'h14)
`define CLP_SHA512_ACC_CSR_EXECUTE                                                                  (32'h30021018)
`define SHA512_ACC_CSR_EXECUTE                                                                      (32'h18)
`define SHA512_ACC_CSR_EXECUTE_EXECUTE_LOW                                                          (0)
`define SHA512_ACC_CSR_EXECUTE_EXECUTE_MASK                                                         (32'h1)
`define CLP_SHA512_ACC_CSR_STATUS                                                                   (32'h3002101c)
`define SHA512_ACC_CSR_STATUS                                                                       (32'h1c)
`define SHA512_ACC_CSR_STATUS_VALID_LOW                                                             (0)
`define SHA512_ACC_CSR_STATUS_VALID_MASK                                                            (32'h1)
`define CLP_SHA512_ACC_CSR_DIGEST_0                                                                 (32'h30021020)
`define SHA512_ACC_CSR_DIGEST_0                                                                     (32'h20)
`define CLP_SHA512_ACC_CSR_DIGEST_1                                                                 (32'h30021024)
`define SHA512_ACC_CSR_DIGEST_1                                                                     (32'h24)
`define CLP_SHA512_ACC_CSR_DIGEST_2                                                                 (32'h30021028)
`define SHA512_ACC_CSR_DIGEST_2                                                                     (32'h28)
`define CLP_SHA512_ACC_CSR_DIGEST_3                                                                 (32'h3002102c)
`define SHA512_ACC_CSR_DIGEST_3                                                                     (32'h2c)
`define CLP_SHA512_ACC_CSR_DIGEST_4                                                                 (32'h30021030)
`define SHA512_ACC_CSR_DIGEST_4                                                                     (32'h30)
`define CLP_SHA512_ACC_CSR_DIGEST_5                                                                 (32'h30021034)
`define SHA512_ACC_CSR_DIGEST_5                                                                     (32'h34)
`define CLP_SHA512_ACC_CSR_DIGEST_6                                                                 (32'h30021038)
`define SHA512_ACC_CSR_DIGEST_6                                                                     (32'h38)
`define CLP_SHA512_ACC_CSR_DIGEST_7                                                                 (32'h3002103c)
`define SHA512_ACC_CSR_DIGEST_7                                                                     (32'h3c)
`define CLP_SHA512_ACC_CSR_DIGEST_8                                                                 (32'h30021040)
`define SHA512_ACC_CSR_DIGEST_8                                                                     (32'h40)
`define CLP_SHA512_ACC_CSR_DIGEST_9                                                                 (32'h30021044)
`define SHA512_ACC_CSR_DIGEST_9                                                                     (32'h44)
`define CLP_SHA512_ACC_CSR_DIGEST_10                                                                (32'h30021048)
`define SHA512_ACC_CSR_DIGEST_10                                                                    (32'h48)
`define CLP_SHA512_ACC_CSR_DIGEST_11                                                                (32'h3002104c)
`define SHA512_ACC_CSR_DIGEST_11                                                                    (32'h4c)
`define CLP_SHA512_ACC_CSR_DIGEST_12                                                                (32'h30021050)
`define SHA512_ACC_CSR_DIGEST_12                                                                    (32'h50)
`define CLP_SHA512_ACC_CSR_DIGEST_13                                                                (32'h30021054)
`define SHA512_ACC_CSR_DIGEST_13                                                                    (32'h54)
`define CLP_SHA512_ACC_CSR_DIGEST_14                                                                (32'h30021058)
`define SHA512_ACC_CSR_DIGEST_14                                                                    (32'h58)
`define CLP_SHA512_ACC_CSR_DIGEST_15                                                                (32'h3002105c)
`define SHA512_ACC_CSR_DIGEST_15                                                                    (32'h5c)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_START                                                      (32'h30021800)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                           (32'h30021800)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h800)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                  (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                 (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                  (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                 (32'h2)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R                                            (32'h30021804)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h804)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                  (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                 (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                  (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                 (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                  (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                 (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                  (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                 (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                            (32'h30021808)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h808)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                          (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                         (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                        (32'h3002180c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h80c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                               (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                        (32'h30021810)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h810)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                               (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                      (32'h30021814)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h814)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                           (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                          (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                           (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                          (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                           (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                          (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                           (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                          (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                      (32'h30021818)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h818)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                   (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                  (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                          (32'h3002181c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h81c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                              (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                             (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                              (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                             (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                              (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                             (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                              (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                             (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                          (32'h30021820)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h820)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                      (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                     (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                        (32'h30021900)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h900)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                        (32'h30021904)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h904)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                        (32'h30021908)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h908)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                        (32'h3002190c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h90c)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                (32'h30021980)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h980)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                   (32'h30021a00)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'ha00)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                   (32'h30021a04)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'ha04)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                   (32'h30021a08)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'ha08)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                   (32'h30021a0c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'ha0c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                           (32'h30021a10)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'ha10)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                     (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                    (32'h1)
`define CLP_SOC_IFC_REG_BASE_ADDR                                                                   (32'h30030000)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_FATAL                                                        (32'h30030000)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL                                                            (32'h0)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL                                                    (32'h30030004)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL                                                        (32'h4)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_FATAL                                                        (32'h30030008)
`define SOC_IFC_REG_CPTRA_FW_ERROR_FATAL                                                            (32'h8)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_NON_FATAL                                                    (32'h3003000c)
`define SOC_IFC_REG_CPTRA_FW_ERROR_NON_FATAL                                                        (32'hc)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_ENC                                                          (32'h30030010)
`define SOC_IFC_REG_CPTRA_HW_ERROR_ENC                                                              (32'h10)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_ENC                                                          (32'h30030014)
`define SOC_IFC_REG_CPTRA_FW_ERROR_ENC                                                              (32'h14)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                              (32'h30030018)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                                  (32'h18)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                              (32'h3003001c)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                                  (32'h1c)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                              (32'h30030020)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                                  (32'h20)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                              (32'h30030024)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                                  (32'h24)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                              (32'h30030028)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                                  (32'h28)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                              (32'h3003002c)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                                  (32'h2c)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                              (32'h30030030)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                                  (32'h30)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                              (32'h30030034)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                                  (32'h34)
`define CLP_SOC_IFC_REG_CPTRA_BOOT_STATUS                                                           (32'h30030038)
`define SOC_IFC_REG_CPTRA_BOOT_STATUS                                                               (32'h38)
`define CLP_SOC_IFC_REG_CPTRA_FLOW_STATUS                                                           (32'h3003003c)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS                                                               (32'h3c)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_STATUS_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_STATUS_MASK                                                   (32'hfffffff)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FW_LOW                                              (28)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FW_MASK                                             (32'h10000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_RUNTIME_LOW                                         (29)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_RUNTIME_MASK                                        (32'h20000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FUSES_LOW                                           (30)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FUSES_MASK                                          (32'h40000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_MAILBOX_FLOW_DONE_LOW                                         (31)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_MAILBOX_FLOW_DONE_MASK                                        (32'h80000000)
`define CLP_SOC_IFC_REG_CPTRA_RESET_REASON                                                          (32'h30030040)
`define SOC_IFC_REG_CPTRA_RESET_REASON                                                              (32'h40)
`define SOC_IFC_REG_CPTRA_RESET_REASON_FW_UPD_RESET_LOW                                             (0)
`define SOC_IFC_REG_CPTRA_RESET_REASON_FW_UPD_RESET_MASK                                            (32'h1)
`define SOC_IFC_REG_CPTRA_RESET_REASON_WARM_RESET_LOW                                               (1)
`define SOC_IFC_REG_CPTRA_RESET_REASON_WARM_RESET_MASK                                              (32'h2)
`define CLP_SOC_IFC_REG_CPTRA_SECURITY_STATE                                                        (32'h30030044)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE                                                            (32'h44)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEVICE_LIFECYCLE_LOW                                       (0)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEVICE_LIFECYCLE_MASK                                      (32'h3)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEBUG_LOCKED_LOW                                           (2)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEBUG_LOCKED_MASK                                          (32'h4)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_RSVD_LOW                                                   (3)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_RSVD_MASK                                                  (32'hfffffff8)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_0                                                        (32'h30030048)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_0                                                            (32'h48)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_1                                                        (32'h3003004c)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_1                                                            (32'h4c)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_2                                                        (32'h30030050)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_2                                                            (32'h50)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_3                                                        (32'h30030054)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_3                                                            (32'h54)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_4                                                        (32'h30030058)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_4                                                            (32'h58)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_0                                                         (32'h3003005c)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_0                                                             (32'h5c)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_0_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_0_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_1                                                         (32'h30030060)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_1                                                             (32'h60)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_1_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_1_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_2                                                         (32'h30030064)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_2                                                             (32'h64)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_2_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_2_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_3                                                         (32'h30030068)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_3                                                             (32'h68)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_3_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_3_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_4                                                         (32'h3003006c)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_4                                                             (32'h6c)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_4_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_4_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_VALID_PAUSER                                                     (32'h30030070)
`define SOC_IFC_REG_CPTRA_TRNG_VALID_PAUSER                                                         (32'h70)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_PAUSER_LOCK                                                      (32'h30030074)
`define SOC_IFC_REG_CPTRA_TRNG_PAUSER_LOCK                                                          (32'h74)
`define SOC_IFC_REG_CPTRA_TRNG_PAUSER_LOCK_LOCK_LOW                                                 (0)
`define SOC_IFC_REG_CPTRA_TRNG_PAUSER_LOCK_LOCK_MASK                                                (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_0                                                           (32'h30030078)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_0                                                               (32'h78)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_1                                                           (32'h3003007c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_1                                                               (32'h7c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_2                                                           (32'h30030080)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_2                                                               (32'h80)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_3                                                           (32'h30030084)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_3                                                               (32'h84)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_4                                                           (32'h30030088)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_4                                                               (32'h88)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_5                                                           (32'h3003008c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_5                                                               (32'h8c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_6                                                           (32'h30030090)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_6                                                               (32'h90)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_7                                                           (32'h30030094)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_7                                                               (32'h94)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_8                                                           (32'h30030098)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_8                                                               (32'h98)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_9                                                           (32'h3003009c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_9                                                               (32'h9c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_10                                                          (32'h300300a0)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_10                                                              (32'ha0)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_11                                                          (32'h300300a4)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_11                                                              (32'ha4)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_STATUS                                                           (32'h300300a8)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS                                                               (32'ha8)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_REQ_LOW                                                  (0)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_REQ_MASK                                                 (32'h1)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_WR_DONE_LOW                                              (1)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_WR_DONE_MASK                                             (32'h2)
`define CLP_SOC_IFC_REG_CPTRA_FUSE_WR_DONE                                                          (32'h300300ac)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE                                                              (32'hac)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE_DONE_LOW                                                     (0)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE_DONE_MASK                                                    (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TIMER_CONFIG                                                          (32'h300300b0)
`define SOC_IFC_REG_CPTRA_TIMER_CONFIG                                                              (32'hb0)
`define CLP_SOC_IFC_REG_CPTRA_BOOTFSM_GO                                                            (32'h300300b4)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO                                                                (32'hb4)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO_GO_LOW                                                         (0)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO_GO_MASK                                                        (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG                                                 (32'h300300b8)
`define SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG                                                     (32'hb8)
`define CLP_SOC_IFC_REG_CPTRA_CLK_GATING_EN                                                         (32'h300300bc)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN                                                             (32'hbc)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN_CLK_GATING_EN_LOW                                           (0)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN_CLK_GATING_EN_MASK                                          (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_0                                                 (32'h300300c0)
`define SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_0                                                     (32'hc0)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_1                                                 (32'h300300c4)
`define SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_1                                                     (32'hc4)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                                (32'h300300c8)
`define SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                                    (32'hc8)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                                (32'h300300cc)
`define SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                                    (32'hcc)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_0                                                             (32'h30030200)
`define SOC_IFC_REG_FUSE_UDS_SEED_0                                                                 (32'h200)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_1                                                             (32'h30030204)
`define SOC_IFC_REG_FUSE_UDS_SEED_1                                                                 (32'h204)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_2                                                             (32'h30030208)
`define SOC_IFC_REG_FUSE_UDS_SEED_2                                                                 (32'h208)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_3                                                             (32'h3003020c)
`define SOC_IFC_REG_FUSE_UDS_SEED_3                                                                 (32'h20c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_4                                                             (32'h30030210)
`define SOC_IFC_REG_FUSE_UDS_SEED_4                                                                 (32'h210)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_5                                                             (32'h30030214)
`define SOC_IFC_REG_FUSE_UDS_SEED_5                                                                 (32'h214)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_6                                                             (32'h30030218)
`define SOC_IFC_REG_FUSE_UDS_SEED_6                                                                 (32'h218)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_7                                                             (32'h3003021c)
`define SOC_IFC_REG_FUSE_UDS_SEED_7                                                                 (32'h21c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_8                                                             (32'h30030220)
`define SOC_IFC_REG_FUSE_UDS_SEED_8                                                                 (32'h220)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_9                                                             (32'h30030224)
`define SOC_IFC_REG_FUSE_UDS_SEED_9                                                                 (32'h224)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_10                                                            (32'h30030228)
`define SOC_IFC_REG_FUSE_UDS_SEED_10                                                                (32'h228)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_11                                                            (32'h3003022c)
`define SOC_IFC_REG_FUSE_UDS_SEED_11                                                                (32'h22c)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_0                                                        (32'h30030230)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_0                                                            (32'h230)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_1                                                        (32'h30030234)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_1                                                            (32'h234)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_2                                                        (32'h30030238)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_2                                                            (32'h238)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_3                                                        (32'h3003023c)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_3                                                            (32'h23c)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_4                                                        (32'h30030240)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_4                                                            (32'h240)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_5                                                        (32'h30030244)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_5                                                            (32'h244)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_6                                                        (32'h30030248)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_6                                                            (32'h248)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_7                                                        (32'h3003024c)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_7                                                            (32'h24c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_0                                                 (32'h30030250)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_0                                                     (32'h250)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_1                                                 (32'h30030254)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_1                                                     (32'h254)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_2                                                 (32'h30030258)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_2                                                     (32'h258)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_3                                                 (32'h3003025c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_3                                                     (32'h25c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_4                                                 (32'h30030260)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_4                                                     (32'h260)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_5                                                 (32'h30030264)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_5                                                     (32'h264)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_6                                                 (32'h30030268)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_6                                                     (32'h268)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_7                                                 (32'h3003026c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_7                                                     (32'h26c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_8                                                 (32'h30030270)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_8                                                     (32'h270)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_9                                                 (32'h30030274)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_9                                                     (32'h274)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_10                                                (32'h30030278)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_10                                                    (32'h278)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_11                                                (32'h3003027c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_11                                                    (32'h27c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK                                              (32'h30030280)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK                                                  (32'h280)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK_MASK_LOW                                         (0)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK_MASK_MASK                                        (32'hf)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_0                                                        (32'h30030284)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_0                                                            (32'h284)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_1                                                        (32'h30030288)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_1                                                            (32'h288)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_2                                                        (32'h3003028c)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_2                                                            (32'h28c)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_3                                                        (32'h30030290)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_3                                                            (32'h290)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_4                                                        (32'h30030294)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_4                                                            (32'h294)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_5                                                        (32'h30030298)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_5                                                            (32'h298)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_6                                                        (32'h3003029c)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_6                                                            (32'h29c)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_7                                                        (32'h300302a0)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_7                                                            (32'h2a0)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_8                                                        (32'h300302a4)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_8                                                            (32'h2a4)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_9                                                        (32'h300302a8)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_9                                                            (32'h2a8)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_10                                                       (32'h300302ac)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_10                                                           (32'h2ac)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_11                                                       (32'h300302b0)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_11                                                           (32'h2b0)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_SVN                                                       (32'h300302b4)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_SVN                                                           (32'h2b4)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_0                                                          (32'h300302b8)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_0                                                              (32'h2b8)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_1                                                          (32'h300302bc)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_1                                                              (32'h2bc)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_2                                                          (32'h300302c0)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_2                                                              (32'h2c0)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_3                                                          (32'h300302c4)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_3                                                              (32'h2c4)
`define CLP_SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE                                                  (32'h300302c8)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE                                                      (32'h2c8)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE_DIS_LOW                                              (0)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE_DIS_MASK                                             (32'h1)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_0                                                     (32'h300302cc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_0                                                         (32'h2cc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_1                                                     (32'h300302d0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_1                                                         (32'h2d0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_2                                                     (32'h300302d4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_2                                                         (32'h2d4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_3                                                     (32'h300302d8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_3                                                         (32'h2d8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_4                                                     (32'h300302dc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_4                                                         (32'h2dc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_5                                                     (32'h300302e0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_5                                                         (32'h2e0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6                                                     (32'h300302e4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6                                                         (32'h2e4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7                                                     (32'h300302e8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7                                                         (32'h2e8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8                                                     (32'h300302ec)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8                                                         (32'h2ec)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9                                                     (32'h300302f0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9                                                         (32'h2f0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10                                                    (32'h300302f4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10                                                        (32'h2f4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_11                                                    (32'h300302f8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_11                                                        (32'h2f8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_12                                                    (32'h300302fc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_12                                                        (32'h2fc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_13                                                    (32'h30030300)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_13                                                        (32'h300)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_14                                                    (32'h30030304)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_14                                                        (32'h304)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_15                                                    (32'h30030308)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_15                                                        (32'h308)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_16                                                    (32'h3003030c)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_16                                                        (32'h30c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_17                                                    (32'h30030310)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_17                                                        (32'h310)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_18                                                    (32'h30030314)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_18                                                        (32'h314)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_19                                                    (32'h30030318)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_19                                                        (32'h318)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_20                                                    (32'h3003031c)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_20                                                        (32'h31c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_21                                                    (32'h30030320)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_21                                                        (32'h320)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_22                                                    (32'h30030324)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_22                                                        (32'h324)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_23                                                    (32'h30030328)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_23                                                        (32'h328)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                                  (32'h3003032c)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                                      (32'h32c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                                  (32'h30030330)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                                      (32'h330)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                                  (32'h30030334)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                                      (32'h334)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                                  (32'h30030338)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                                      (32'h338)
`define CLP_SOC_IFC_REG_FUSE_LIFE_CYCLE                                                             (32'h3003033c)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE                                                                 (32'h33c)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE_LIFE_CYCLE_LOW                                                  (0)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE_LIFE_CYCLE_MASK                                                 (32'h3)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_0                                                          (32'h30030600)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_0                                                              (32'h600)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_1                                                          (32'h30030604)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_1                                                              (32'h604)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_2                                                          (32'h30030608)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_2                                                              (32'h608)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_3                                                          (32'h3003060c)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_3                                                              (32'h60c)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_4                                                          (32'h30030610)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_4                                                              (32'h610)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_5                                                          (32'h30030614)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_5                                                              (32'h614)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_6                                                          (32'h30030618)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_6                                                              (32'h618)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_7                                                          (32'h3003061c)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_7                                                              (32'h61c)
`define CLP_SOC_IFC_REG_INTERNAL_ICCM_LOCK                                                          (32'h30030620)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK                                                              (32'h620)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK_LOCK_LOW                                                     (0)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK_LOCK_MASK                                                    (32'h1)
`define CLP_SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET                                                    (32'h30030624)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET                                                        (32'h624)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_CORE_RST_LOW                                           (0)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_CORE_RST_MASK                                          (32'h1)
`define CLP_SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES                                        (32'h30030628)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES                                            (32'h628)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES_WAIT_CYCLES_LOW                            (0)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES_WAIT_CYCLES_MASK                           (32'hff)
`define CLP_SOC_IFC_REG_INTERNAL_NMI_VECTOR                                                         (32'h3003062c)
`define SOC_IFC_REG_INTERNAL_NMI_VECTOR                                                             (32'h62c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_START                                                         (32'h30030800)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                              (32'h30030800)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h800)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                     (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                    (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                     (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                    (32'h2)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                               (32'h30030804)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h804)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_LOW                             (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_MASK                            (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INV_DEV_EN_LOW                              (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INV_DEV_EN_MASK                             (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_CMD_FAIL_EN_LOW                             (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_CMD_FAIL_EN_MASK                            (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_BAD_FUSE_EN_LOW                             (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_BAD_FUSE_EN_MASK                            (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_ICCM_BLOCKED_EN_LOW                         (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_ICCM_BLOCKED_EN_MASK                        (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_MBOX_ECC_UNC_EN_LOW                         (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_MBOX_ECC_UNC_EN_MASK                        (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                               (32'h30030808)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h808)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_AVAIL_EN_LOW                            (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_AVAIL_EN_MASK                           (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_MBOX_ECC_COR_EN_LOW                         (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_MBOX_ECC_COR_EN_MASK                        (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_DEBUG_LOCKED_EN_LOW                         (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_DEBUG_LOCKED_EN_MASK                        (32'h4)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                           (32'h3003080c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h80c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                   (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                  (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                           (32'h30030810)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h810)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                   (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                  (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                         (32'h30030814)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h814)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_LOW                      (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_MASK                     (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INV_DEV_STS_LOW                       (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INV_DEV_STS_MASK                      (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_CMD_FAIL_STS_LOW                      (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_CMD_FAIL_STS_MASK                     (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_BAD_FUSE_STS_LOW                      (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_BAD_FUSE_STS_MASK                     (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_ICCM_BLOCKED_STS_LOW                  (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_ICCM_BLOCKED_STS_MASK                 (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_MBOX_ECC_UNC_STS_LOW                  (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_MBOX_ECC_UNC_STS_MASK                 (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                         (32'h30030818)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h818)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_AVAIL_STS_LOW                     (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_AVAIL_STS_MASK                    (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_MBOX_ECC_COR_STS_LOW                  (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_MBOX_ECC_COR_STS_MASK                 (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_DEBUG_LOCKED_STS_LOW                  (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_DEBUG_LOCKED_STS_MASK                 (32'h4)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                             (32'h3003081c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h81c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_LOW                         (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_MASK                        (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INV_DEV_TRIG_LOW                          (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INV_DEV_TRIG_MASK                         (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_CMD_FAIL_TRIG_LOW                         (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_CMD_FAIL_TRIG_MASK                        (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_BAD_FUSE_TRIG_LOW                         (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_BAD_FUSE_TRIG_MASK                        (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_ICCM_BLOCKED_TRIG_LOW                     (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_ICCM_BLOCKED_TRIG_MASK                    (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_MBOX_ECC_UNC_TRIG_LOW                     (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_MBOX_ECC_UNC_TRIG_MASK                    (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                             (32'h30030820)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h820)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_AVAIL_TRIG_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_AVAIL_TRIG_MASK                       (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_MBOX_ECC_COR_TRIG_LOW                     (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_MBOX_ECC_COR_TRIG_MASK                    (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_DEBUG_LOCKED_TRIG_LOW                     (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_DEBUG_LOCKED_TRIG_MASK                    (32'h4)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                   (32'h30030900)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h900)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_R                                    (32'h30030904)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_R                                        (32'h904)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_R                                   (32'h30030908)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_R                                       (32'h908)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_R                                   (32'h3003090c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_R                                       (32'h90c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_R                               (32'h30030910)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_R                                   (32'h910)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_R                               (32'h30030914)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_R                                   (32'h914)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_R                                  (32'h30030980)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_R                                      (32'h980)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_R                               (32'h30030984)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_R                                   (32'h984)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                               (32'h30030988)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                                   (32'h988)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                              (32'h30030a00)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'ha00)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R                               (32'h30030a04)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R                                   (32'ha04)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R                              (32'h30030a08)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R                                  (32'ha08)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R                              (32'h30030a0c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R                                  (32'ha0c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R                          (32'h30030a10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R                              (32'ha10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R                          (32'h30030a14)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R                              (32'ha14)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R                             (32'h30030a18)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R                                 (32'ha18)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R_PULSE_LOW                       (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R_PULSE_MASK                      (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R                          (32'h30030a1c)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R                              (32'ha1c)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                          (32'h30030a20)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                              (32'ha20)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)


`endif