//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This interface performs the pv_write signal monitoring.
//      It is accessed by the uvm pv_write monitor through a virtual
//      interface handle in the pv_write configuration.  It monitors the
//      signals passed in through the port connection named bus of
//      type pv_write_if.
//
//     Input signals from the pv_write_if are assigned to an internal input
//     signal with a _i suffix.  The _i signal should be used for sampling.
//
//     The input signal connections are as follows:
//       bus.signal -> signal_i 
//
//      Interface functions and tasks used by UVM components:
//             monitor(inout TRANS_T txn);
//                   This task receives the transaction, txn, from the
//                   UVM monitor and then populates variables in txn
//                   from values observed on bus activity.  This task
//                   blocks until an operation on the pv_write bus is complete.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
import uvmf_base_pkg_hdl::*;
import pv_write_pkg_hdl::*;
`include "src/pv_write_macros.svh"


interface pv_write_monitor_bfm #(
  string PV_WRITE_REQUESTOR = "SHA512"
  )

  ( pv_write_if  bus );
  // The pragma below and additional ones in-lined further down are for running this BFM on Veloce
  // pragma attribute pv_write_monitor_bfm partition_interface_xif                                  

`ifndef XRTL
// This code is to aid in debugging parameter mismatches between the BFM and its corresponding agent.
// Enable this debug by setting UVM_VERBOSITY to UVM_DEBUG
// Setting UVM_VERBOSITY to UVM_DEBUG causes all BFM's and all agents to display their parameter settings.
// All of the messages from this feature have a UVM messaging id value of "CFG"
// The transcript or run.log can be parsed to ensure BFM parameter settings match its corresponding agents parameter settings.
import uvm_pkg::*;
`include "uvm_macros.svh"
initial begin : bfm_vs_agent_parameter_debug
  `uvm_info("CFG", 
      $psprintf("The BFM at '%m' has the following parameters: PV_WRITE_REQUESTOR=%x ", PV_WRITE_REQUESTOR),
      UVM_DEBUG)
end
`endif


  // Structure used to pass transaction data from monitor BFM to monitor class in agent.
`pv_write_MONITOR_STRUCT
  pv_write_monitor_s pv_write_monitor_struct;

  // Structure used to pass configuration data from monitor class to monitor BFM.
 `pv_write_CONFIGURATION_STRUCT
 

  // Config value to determine if this is an initiator or a responder 
  uvmf_initiator_responder_t initiator_responder;
  // Custom configuration variables.  
  // These are set using the configure function which is called during the UVM connect_phase

  tri clk_i;
  tri dummy_i;
  tri [$bits(pv_defines_pkg::pv_write_t)-1:0] pv_write_i;
  tri [$bits(pv_defines_pkg::pv_wr_resp_t)-1:0] pv_wr_resp_i;

  reg write_en_i;
  reg [PV_ENTRY_ADDR_W-1:0] write_entry_i;
  reg [PV_ENTRY_SIZE_WIDTH-1:0] write_offset_i;
  reg [PV_DATA_W-1:0] write_data_i;
  reg error_i;

  assign clk_i = bus.clk;
  assign dummy_i = bus.dummy;
  assign pv_write_i = bus.pv_write;
  assign pv_wr_resp_i = bus.pv_wr_resp;

  assign write_en_i          = pv_write_i[41]; 
  assign write_entry_i       = pv_write_i[40:36]; 
  assign write_offset_i      = pv_write_i[35:32]; 
  assign write_data_i        = pv_write_i[31:0]; 

  assign error_i             = pv_wr_resp_i[0];

  // Proxy handle to UVM monitor
  pv_write_pkg::pv_write_monitor #(
    .PV_WRITE_REQUESTOR(PV_WRITE_REQUESTOR)
    )
 proxy;
  // pragma tbx oneway proxy.notify_transaction                 

  // pragma uvmf custom interface_item_additional begin
 reg write_en_o                               = 'h0; 
 reg [PV_ENTRY_ADDR_W-1:0] write_entry_o      = 'h0; 
 reg [PV_ENTRY_SIZE_WIDTH-1:0] write_offset_o     = 'h0; 
 reg [PV_DATA_W-1:0] write_data_o             = 'h0; 
 
 reg error_o = 'h0;

 function any_signal_changed();

  return |(write_en_i ^ write_en_o) ||
         |(write_entry_i ^ write_entry_o) ||
         |(write_offset_i ^ write_offset_o) ||
         |(write_data_i ^ write_data_o) ; //||
         //|(error_i ^ error_o);

 endfunction
  // pragma uvmf custom interface_item_additional end
  
  //******************************************************************                         
  task wait_for_reset();// pragma tbx xtf  
    @(posedge clk_i) ;                                                                    
    do_wait_for_reset();                                                                   
  endtask                                                                                   

  // ****************************************************************************              
  task do_wait_for_reset(); 
  // pragma uvmf custom reset_condition begin
    wait ( dummy_i === 1 ) ;                                                              
    @(posedge clk_i) ;                                                                    
  // pragma uvmf custom reset_condition end                                                                
  endtask    

  //******************************************************************                         
 
  task wait_for_num_clocks(input int unsigned count); // pragma tbx xtf 
    @(posedge clk_i);  
                                                                   
    repeat (count-1) @(posedge clk_i);                                                    
  endtask      

  //******************************************************************                         
  event go;                                                                                 
  function void start_monitoring();// pragma tbx xtf    
    -> go;
  endfunction                                                                               
  
  // ****************************************************************************              
  initial begin                                                                             
    @go;                                                                                   
    forever begin                                                                        
      //@(posedge clk_i);  //No delay between DRV and MON to make sure PRED receives txn in time
      do_monitor( pv_write_monitor_struct );
                                                                 
 
      proxy.notify_transaction( pv_write_monitor_struct );
 
    end                                                                                    
  end                                                                                       

  //******************************************************************
  // The configure() function is used to pass agent configuration
  // variables to the monitor BFM.  It is called by the monitor within
  // the agent at the beginning of the simulation.  It may be called 
  // during the simulation if agent configuration variables are updated
  // and the monitor BFM needs to be aware of the new configuration 
  // variables.
  //
    function void configure(pv_write_configuration_s pv_write_configuration_arg); // pragma tbx xtf  
    initiator_responder = pv_write_configuration_arg.initiator_responder;
  // pragma uvmf custom configure begin
  // pragma uvmf custom configure end
  endfunction   


  // ****************************************************************************  
            
  task do_monitor(output pv_write_monitor_s pv_write_monitor_struct);
    //
    // Available struct members:
    //     //    pv_write_monitor_struct.write_en
    //     //    pv_write_monitor_struct.write_entry
    //     //    pv_write_monitor_struct.write_offset
    //     //    pv_write_monitor_struct.write_data
    //     //    pv_write_monitor_struct.error
    //     //
    // Reference code;
    //    How to wait for signal value
    //      while (control_signal === 1'b1) @(posedge clk_i);
    //    
    //    How to assign a struct member, named xyz, from a signal.   
    //    All available input signals listed.
    //      pv_write_monitor_struct.xyz = pv_write_i;  //    [$bits(pv_defines_pkg::pv_write_t)-1:0] 
    //      pv_write_monitor_struct.xyz = pv_wr_resp_i;  //    [$bits(pv_defines_pkg::pv_wr_resp_t)-1:0] 
    // pragma uvmf custom do_monitor begin
    // UVMF_CHANGE_ME : Implement protocol monitoring.  The commented reference code 
    // below are examples of how to capture signal values and assign them to 
    // structure members.  All available input signals are listed.  The 'while' 
    // code example shows how to wait for a synchronous flow control signal.  This
    // task should return when a complete transfer has been observed.  Once this task is
    // exited with captured values, it is then called again to wait for and observe 
    // the next transfer. One clock cycle is consumed between calls to do_monitor.
    while(!any_signal_changed()) @(posedge clk_i);
    write_en_o          <= write_en_i;
    write_entry_o       <= write_entry_i;
    write_offset_o      <= write_offset_i;
    write_data_o        <= write_data_i;
    error_o             <= error_i;

    @(posedge clk_i); //Delay write txn to monitor by 1 clk to mimic design
    //(regs are updated in the next clk and reg model should follow the same)

    pv_write_monitor_struct.write_en          = write_en_o;
    pv_write_monitor_struct.write_entry       = write_entry_o;
    pv_write_monitor_struct.write_offset      = write_offset_o;
    pv_write_monitor_struct.write_data        = write_data_o;
    pv_write_monitor_struct.error             = error_o;

    // pragma uvmf custom do_monitor end
  endtask         
  
 
endinterface

// pragma uvmf custom external begin
// pragma uvmf custom external end

