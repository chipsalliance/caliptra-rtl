  //----------------------------------------------------------------
  // Internal constant and parameter definitions.
  //----------------------------------------------------------------
  localparam HMAC_DRBG_SEED_LENGTH        = 32'd384;
  