// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef CALIPTRA_TOP_REG_DEFINES_HEADER
`define CALIPTRA_TOP_REG_DEFINES_HEADER


`define CALIPTRA_TOP_REG_BASE_ADDR                                                                  (32'h0)
`define CALIPTRA_TOP_REG_MBOX_CSR_BASE_ADDR                                                         (32'h20000)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_LOCK                                                         (32'h20000)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_USER                                                         (32'h20004)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_CMD                                                          (32'h20008)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_DLEN                                                         (32'h2000c)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_DATAIN                                                       (32'h20010)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_DATAOUT                                                      (32'h20014)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_EXECUTE                                                      (32'h20018)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_STATUS                                                       (32'h2001c)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_UNLOCK                                                       (32'h20020)
`define CALIPTRA_TOP_REG_MBOX_CSR_TAP_MODE                                                          (32'h20024)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_BASE_ADDR                                             (32'h30000)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL                                  (32'h30000)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL                              (32'h30004)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_FATAL                                  (32'h30008)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_NON_FATAL                              (32'h3000c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_ENC                                    (32'h30010)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_ENC                                    (32'h30014)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                        (32'h30018)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                        (32'h3001c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                        (32'h30020)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                        (32'h30024)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                        (32'h30028)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                        (32'h3002c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                        (32'h30030)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                        (32'h30034)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_BOOT_STATUS                                     (32'h30038)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS                                     (32'h3003c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_RESET_REASON                                    (32'h30040)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE                                  (32'h30044)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_AXI_USER_0                           (32'h30048)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_AXI_USER_1                           (32'h3004c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_AXI_USER_2                           (32'h30050)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_AXI_USER_3                           (32'h30054)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_AXI_USER_4                           (32'h30058)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_AXI_USER_LOCK_0                            (32'h3005c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_AXI_USER_LOCK_1                            (32'h30060)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_AXI_USER_LOCK_2                            (32'h30064)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_AXI_USER_LOCK_3                            (32'h30068)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_AXI_USER_LOCK_4                            (32'h3006c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_VALID_AXI_USER                             (32'h30070)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_AXI_USER_LOCK                              (32'h30074)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_0                                     (32'h30078)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_1                                     (32'h3007c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_2                                     (32'h30080)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_3                                     (32'h30084)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_4                                     (32'h30088)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_5                                     (32'h3008c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_6                                     (32'h30090)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_7                                     (32'h30094)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_8                                     (32'h30098)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_9                                     (32'h3009c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_10                                    (32'h300a0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_11                                    (32'h300a4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_CTRL                                       (32'h300a8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_STATUS                                     (32'h300ac)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FUSE_WR_DONE                                    (32'h300b0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TIMER_CONFIG                                    (32'h300b4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_BOOTFSM_GO                                      (32'h300b8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_DBG_MANUF_SERVICE_REG                           (32'h300bc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_CLK_GATING_EN                                   (32'h300c0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_GENERIC_INPUT_WIRES_0                           (32'h300c4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_GENERIC_INPUT_WIRES_1                           (32'h300c8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                          (32'h300cc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                          (32'h300d0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_REV_ID                                       (32'h300d4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_REV_ID_0                                     (32'h300d8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_REV_ID_1                                     (32'h300dc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG                                       (32'h300e0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_EN                                   (32'h300e4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_CTRL                                 (32'h300e8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_0                     (32'h300ec)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_1                     (32'h300f0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_EN                                   (32'h300f4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_CTRL                                 (32'h300f8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_0                     (32'h300fc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_1                     (32'h30100)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_STATUS                                      (32'h30104)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FUSE_VALID_AXI_USER                             (32'h30108)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FUSE_AXI_USER_LOCK                              (32'h3010c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_CFG_0                                       (32'h30110)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_CFG_1                                       (32'h30114)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0                          (32'h30118)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1                          (32'h3011c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_RSVD_REG_0                                      (32'h30120)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_RSVD_REG_1                                      (32'h30124)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_CAPABILITIES                                 (32'h30128)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_CAPABILITIES                                 (32'h3012c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_CAP_LOCK                                        (32'h30130)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_0                                 (32'h30140)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_1                                 (32'h30144)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_2                                 (32'h30148)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_3                                 (32'h3014c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_4                                 (32'h30150)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_5                                 (32'h30154)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_6                                 (32'h30158)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_7                                 (32'h3015c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_8                                 (32'h30160)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_9                                 (32'h30164)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_10                                (32'h30168)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_11                                (32'h3016c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_OWNER_PK_HASH_LOCK                              (32'h30170)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_0                                       (32'h30200)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_1                                       (32'h30204)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_2                                       (32'h30208)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_3                                       (32'h3020c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_4                                       (32'h30210)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_5                                       (32'h30214)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_6                                       (32'h30218)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_7                                       (32'h3021c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_8                                       (32'h30220)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_9                                       (32'h30224)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_10                                      (32'h30228)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_11                                      (32'h3022c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_12                                      (32'h30230)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_13                                      (32'h30234)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_14                                      (32'h30238)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_15                                      (32'h3023c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_0                                  (32'h30240)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_1                                  (32'h30244)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_2                                  (32'h30248)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_3                                  (32'h3024c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_4                                  (32'h30250)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_5                                  (32'h30254)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_6                                  (32'h30258)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_7                                  (32'h3025c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_0                                 (32'h30260)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_1                                 (32'h30264)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_2                                 (32'h30268)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_3                                 (32'h3026c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_4                                 (32'h30270)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_5                                 (32'h30274)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_6                                 (32'h30278)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_7                                 (32'h3027c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_8                                 (32'h30280)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_9                                 (32'h30284)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_10                                (32'h30288)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_VENDOR_PK_HASH_11                                (32'h3028c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_ECC_REVOCATION                                   (32'h30290)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FMC_KEY_MANIFEST_SVN                             (32'h302b4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_0                                    (32'h302b8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_1                                    (32'h302bc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_2                                    (32'h302c0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_3                                    (32'h302c4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_ANTI_ROLLBACK_DISABLE                            (32'h302c8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_0                               (32'h302cc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_1                               (32'h302d0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_2                               (32'h302d4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_3                               (32'h302d8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_4                               (32'h302dc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_5                               (32'h302e0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_6                               (32'h302e4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_7                               (32'h302e8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_8                               (32'h302ec)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_9                               (32'h302f0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_10                              (32'h302f4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_11                              (32'h302f8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_12                              (32'h302fc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_13                              (32'h30300)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_14                              (32'h30304)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_15                              (32'h30308)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_16                              (32'h3030c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_17                              (32'h30310)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_18                              (32'h30314)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_19                              (32'h30318)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_20                              (32'h3031c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_21                              (32'h30320)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_22                              (32'h30324)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_23                              (32'h30328)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_0                            (32'h3032c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_1                            (32'h30330)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_2                            (32'h30334)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_3                            (32'h30338)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_LMS_REVOCATION                                   (32'h30340)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_MLDSA_REVOCATION                                 (32'h30344)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_SOC_STEPPING_ID                                  (32'h30348)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_0                         (32'h3034c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_1                         (32'h30350)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_2                         (32'h30354)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_3                         (32'h30358)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_PQC_KEY_TYPE                                     (32'h3035c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_SOC_MANIFEST_SVN_0                               (32'h30360)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_SOC_MANIFEST_SVN_1                               (32'h30364)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_SOC_MANIFEST_SVN_2                               (32'h30368)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_SOC_MANIFEST_SVN_3                               (32'h3036c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_SOC_MANIFEST_MAX_SVN                             (32'h30370)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_CALIPTRA_BASE_ADDR_L                               (32'h30500)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_CALIPTRA_BASE_ADDR_H                               (32'h30504)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_MCI_BASE_ADDR_L                                    (32'h30508)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_MCI_BASE_ADDR_H                                    (32'h3050c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_RECOVERY_IFC_BASE_ADDR_L                           (32'h30510)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_RECOVERY_IFC_BASE_ADDR_H                           (32'h30514)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_OTP_FC_BASE_ADDR_L                                 (32'h30518)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_OTP_FC_BASE_ADDR_H                                 (32'h3051c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_UDS_SEED_BASE_ADDR_L                               (32'h30520)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_UDS_SEED_BASE_ADDR_H                               (32'h30524)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_PROD_DEBUG_UNLOCK_AUTH_PK_HASH_REG_BANK_OFFSET     (32'h30528)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_NUM_OF_PROD_DEBUG_UNLOCK_AUTH_PK_HASHES            (32'h3052c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_DEBUG_INTENT                                       (32'h30530)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_CALIPTRA_DMA_AXI_USER                              (32'h30534)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_STRAP_GENERIC_0                                    (32'h305a0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_STRAP_GENERIC_1                                    (32'h305a4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_STRAP_GENERIC_2                                    (32'h305a8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_STRAP_GENERIC_3                                    (32'h305ac)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_DBG_MANUF_SERVICE_REG_REQ                          (32'h305c0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_DBG_MANUF_SERVICE_REG_RSP                          (32'h305c4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_SOC_DBG_UNLOCK_LEVEL_0                             (32'h305c8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_SOC_DBG_UNLOCK_LEVEL_1                             (32'h305cc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_GENERIC_FW_EXEC_CTRL_0                             (32'h305d0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_GENERIC_FW_EXEC_CTRL_1                             (32'h305d4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_GENERIC_FW_EXEC_CTRL_2                             (32'h305d8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_SS_GENERIC_FW_EXEC_CTRL_3                             (32'h305dc)


`endif