// Copyright (C) Microsoft Corporation. All rights reserved.

module integration_tb();
    integration_top integration();
endmodule : integration_tb
