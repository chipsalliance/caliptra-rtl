//
// File: qvip_apb5_slave_pkg.sv
//
// Generated from Mentor VIP Configurator (20220406)
// Generated using Mentor VIP Library ( 2022.2 : 04/20/2022:16:06 )
//
package qvip_apb5_slave_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    import addr_map_pkg::*;
    
    import qvip_apb5_slave_params_pkg::*;
    import mvc_pkg::*;
    import mgc_apb3_v1_0_pkg::*;
    
    `include "qvip_apb5_slave_env_config.svh"
    `include "qvip_apb5_slave_env.svh"
    `include "qvip_apb5_slave_vseq_base.svh"
    `include "qvip_apb5_slave_test_base.svh"
endpackage: qvip_apb5_slave_pkg
