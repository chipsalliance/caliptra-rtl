//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20220406)
// Generated using Mentor VIP Library ( 2022.2 : 04/20/2022:16:06 )
//

import qvip_ahb_lite_slave_test_pkg::*;

// Add other packages here as required
