// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng top level wrapper file

`include "caliptra_prim_assert.sv"

module csrng
 import csrng_pkg::*;
 import csrng_reg_pkg::*;
 import lc_ctrl_state_pkg::*;
 import lc_ctrl_reg_pkg::*;
 import lc_ctrl_pkg::*;
#(
  parameter aes_pkg::sbox_impl_e SBoxImpl = aes_pkg::SBoxImplCanright,
  parameter logic [csrng_reg_pkg::NumAlerts-1:0] AlertAsyncOn = {csrng_reg_pkg::NumAlerts{1'b1}},
  parameter logic [31:0] NHwApps = 2,
  parameter cs_keymgr_div_t RndCnstCsKeymgrDivNonProduction = CsKeymgrDivWidth'(0),
  parameter cs_keymgr_div_t RndCnstCsKeymgrDivProduction = CsKeymgrDivWidth'(0),
  parameter AHBDataWidth = 64,
  parameter AHBAddrWidth = 32
) (
  input logic         clk_i,
  input logic         rst_ni,

  // AMBA AHB Lite Interface
  input logic [AHBAddrWidth-1:0]  haddr_i,
  input logic [AHBDataWidth-1:0]  hwdata_i,
  input logic                     hsel_i,
  input logic                     hwrite_i,
  input logic                     hready_i,
  input logic [1:0]               htrans_i,
  input logic [2:0]               hsize_i,

  output logic                    hresp_o,
  output logic                    hreadyout_o,
  output logic [AHBDataWidth-1:0] hrdata_o,



   // OTP Interface
  // SEC_CM: INTERSIG.MUBI
  input  caliptra_prim_mubi_pkg::mubi8_t otp_en_csrng_sw_app_read_i,

  // Lifecycle broadcast inputs
  input  lc_ctrl_pkg::lc_tx_t  lc_hw_debug_en_i,

  // Entropy Interface
  output entropy_src_pkg::entropy_src_hw_if_req_t entropy_src_hw_if_o,
  input  entropy_src_pkg::entropy_src_hw_if_rsp_t entropy_src_hw_if_i,

  // Entropy Interface
  input  entropy_src_pkg::cs_aes_halt_req_t cs_aes_halt_i,
  output entropy_src_pkg::cs_aes_halt_rsp_t cs_aes_halt_o,

  // Application Interfaces
  input  csrng_req_t  [NHwApps-1:0] csrng_cmd_i,
  output csrng_rsp_t  [NHwApps-1:0] csrng_cmd_o,

  // Alerts
  input  caliptra_prim_alert_pkg::alert_rx_t [csrng_reg_pkg::NumAlerts-1:0] alert_rx_i,
  output caliptra_prim_alert_pkg::alert_tx_t [csrng_reg_pkg::NumAlerts-1:0] alert_tx_o,

  // Interrupts
  output logic    intr_cs_cmd_req_done_o,
  output logic    intr_cs_entropy_req_o,
  output logic    intr_cs_hw_inst_exc_o,
  output logic    intr_cs_fatal_err_o
);

  csrng_reg2hw_t reg2hw;
  csrng_hw2reg_t hw2reg;

  logic [csrng_reg_pkg::NumAlerts-1:0] alert_test;
  logic [csrng_reg_pkg::NumAlerts-1:0] alert;

  logic [csrng_reg_pkg::NumAlerts-1:0] intg_err_alert;
  assign intg_err_alert[0] = 1'b0;

  // SEC_CM: CONFIG.REGWEN
  // SEC_CM: TILE_LINK.BUS.INTEGRITY

  csrng_reg_top #(
    .AHBDataWidth(AHBDataWidth),
    .AHBAddrWidth(AHBAddrWidth)
  ) u_reg (
    .clk_i,
    .rst_ni,
    .haddr_i,
    .hwdata_i,
    .hsel_i,
    .hwrite_i,
    .hready_i,
    .htrans_i,
    .hsize_i,
    .hresp_o,
    .hreadyout_o,
    .hrdata_o,
    .reg2hw,
    .hw2reg,
    .intg_err_o(intg_err_alert[1]),
    .devmode_i(1'b1)
  );

  csrng_core #(
    .SBoxImpl(SBoxImpl),
    .NHwApps(NHwApps),
    .RndCnstCsKeymgrDivNonProduction(RndCnstCsKeymgrDivNonProduction),
    .RndCnstCsKeymgrDivProduction(RndCnstCsKeymgrDivProduction)
  ) u_csrng_core (
    .clk_i,
    .rst_ni,
    .reg2hw,
    .hw2reg,

    // misc inputs
    .otp_en_csrng_sw_app_read_i(otp_en_csrng_sw_app_read_i),
    .lc_hw_debug_en_i,

    // Entropy Interface
    .entropy_src_hw_if_o,
    .entropy_src_hw_if_i,

    // Entropy Interface
    .cs_aes_halt_i,
    .cs_aes_halt_o,

    // Application Interfaces
    .csrng_cmd_i,
    .csrng_cmd_o,

    // Alerts
    .recov_alert_test_o(alert_test[0]),
    .fatal_alert_test_o(alert_test[1]),
    .recov_alert_o(alert[0]),
    .fatal_alert_o(alert[1]),

    .intr_cs_cmd_req_done_o,
    .intr_cs_entropy_req_o,
    .intr_cs_hw_inst_exc_o,
    .intr_cs_fatal_err_o
  );


  ///////////////////////////
  // Alert generation
  ///////////////////////////
  for (genvar i = 0; i < csrng_reg_pkg::NumAlerts; i++) begin : gen_alert_tx
    caliptra_prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(i)
    ) u_caliptra_prim_alert_sender (
      .clk_i,
      .rst_ni,
      .alert_test_i  (alert_test[i]                 ),
      .alert_req_i   (alert[i] || intg_err_alert[i] ),
      .alert_ack_o   (),
      .alert_state_o (),
      .alert_rx_i    (alert_rx_i[i]                 ),
      .alert_tx_o    (alert_tx_o[i]                 )
    );
  end


  // Assertions

  `CALIPTRA_ASSERT_KNOWN(AHBRespKnownO_A, hresp_o)
  `CALIPTRA_ASSERT_KNOWN(AHBReadyKnownO_A, hreadyout_o)
  `CALIPTRA_ASSERT_KNOWN(EsReqKnownO_A, entropy_src_hw_if_o.es_req)

  // Application Interface Asserts
  for (genvar i = 0; i < NHwApps; i = i+1) begin : gen_app_if_asserts
    `CALIPTRA_ASSERT_KNOWN(CsrngReqReadyKnownO_A, csrng_cmd_o[i].csrng_req_ready)
    `CALIPTRA_ASSERT_KNOWN(CsrngRspAckKnownO_A, csrng_cmd_o[i].csrng_rsp_ack)
    `CALIPTRA_ASSERT_KNOWN(CsrngRspStsKnownO_A, csrng_cmd_o[i].csrng_rsp_sts)
    `CALIPTRA_ASSERT_KNOWN(CsrngGenbitsValidKnownO_A, csrng_cmd_o[i].genbits_valid)
    `CALIPTRA_ASSERT_KNOWN(CsrngGenbitsFipsKnownO_A, csrng_cmd_o[i].genbits_fips)
    `CALIPTRA_ASSERT_KNOWN(CsrngGenbitsBusKnownO_A, csrng_cmd_o[i].genbits_bus)
  end : gen_app_if_asserts

  // Alerts
  `CALIPTRA_ASSERT_KNOWN(AlertTxKnownO_A, alert_tx_o)

  `CALIPTRA_ASSERT_KNOWN(IntrCsCmdReqDoneKnownO_A, intr_cs_cmd_req_done_o)
  `CALIPTRA_ASSERT_KNOWN(IntrCsEntropyReqKnownO_A, intr_cs_entropy_req_o)
  `CALIPTRA_ASSERT_KNOWN(IntrCsHwInstExcKnownO_A, intr_cs_hw_inst_exc_o)
  `CALIPTRA_ASSERT_KNOWN(IntrCsFatalErrKnownO_A, intr_cs_fatal_err_o)

  `CALIPTRA_ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CtrDrbgUpdAlertCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_upd.u_caliptra_prim_count_ctr_drbg,
    alert_tx_o[1])

  `CALIPTRA_ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CtrDrbgGenAlertCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_gen.u_caliptra_prim_count_ctr_drbg,
    alert_tx_o[1])

  for (genvar i = 0; i < NHwApps + 1; i++) begin : gen_cnt_asserts
    `CALIPTRA_ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck_A,
      u_csrng_core.gen_cmd_stage[i].u_csrng_cmd_stage.u_caliptra_prim_count_cmd_gen_cntr,
      alert_tx_o[1])

    `CALIPTRA_ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(DrbgCmdFsmCheck_A,
      u_csrng_core.gen_cmd_stage[i].u_csrng_cmd_stage.u_state_regs,
      alert_tx_o[1])
  end

  `CALIPTRA_ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CtrlMainFsmCheck_A,
    u_csrng_core.u_csrng_main_sm.u_state_regs,
    alert_tx_o[1])

  `CALIPTRA_ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(DrbgGenFsmCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_gen.u_state_regs,
    alert_tx_o[1])

  `CALIPTRA_ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(DrbgUpdBlkEncFsmCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_upd.u_blk_enc_state_regs,
    alert_tx_o[1])

  `CALIPTRA_ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(DrbgUpdOutBlkFsmCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_upd.u_outblk_state_regs,
    alert_tx_o[1])

  for (genvar i = 0; i < aes_pkg::Sp2VWidth; i++) begin : gen_aes_cipher_control_fsm_svas
    if (aes_pkg::SP2V_LOGIC_HIGH[i] == 1'b1) begin : gen_aes_cipher_control_fsm_svas_p
      `CALIPTRA_ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesCipherControlFsmCheck_A,
          u_csrng_core.u_csrng_block_encrypt.u_aes_cipher_core.u_aes_cipher_control.gen_fsm[i].
              gen_fsm_p.u_aes_cipher_control_fsm_i.u_aes_cipher_control_fsm.u_state_regs,
          alert_tx_o[1])
    end else begin : gen_aes_cipher_control_fsm_svas_n
      `CALIPTRA_ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesCipherControlFsmCheck_A,
          u_csrng_core.u_csrng_block_encrypt.u_aes_cipher_core.u_aes_cipher_control.gen_fsm[i].
              gen_fsm_n.u_aes_cipher_control_fsm_i.u_aes_cipher_control_fsm.u_state_regs,
          alert_tx_o[1])
    end
  end

  // Alert assertions for reg_we onehot check
  `CALIPTRA_ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A, u_reg, alert_tx_o[1])
endmodule
