//======================================================================
//
// hmac_drbg_tb.sv
//
//
// Author: Emre Karabulut
// 
// This test to check HMAC DRBG functionality
// Empty test
//======================================================================

module hmac_drbg_tb();

endmodule // hmac_drbg_tb

//======================================================================
// EOF hmac_drbg_tb.sv
//======================================================================
