// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef CALIPTRA_TOP_REG_DEFINES_HEADER
`define CALIPTRA_TOP_REG_DEFINES_HEADER


`define CALIPTRA_TOP_REG_BASE_ADDR                                                                  (32'h0)
`define CALIPTRA_TOP_REG_MBOX_CSR_BASE_ADDR                                                         (32'h30020000)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_LOCK                                                         (32'h30020000)
`define MBOX_CSR_MBOX_LOCK                                                                          (32'h0)
`define MBOX_CSR_MBOX_LOCK_LOCK_LOW                                                                 (0)
`define MBOX_CSR_MBOX_LOCK_LOCK_MASK                                                                (32'h1)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_USER                                                         (32'h30020004)
`define MBOX_CSR_MBOX_USER                                                                          (32'h4)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_CMD                                                          (32'h30020008)
`define MBOX_CSR_MBOX_CMD                                                                           (32'h8)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_DLEN                                                         (32'h3002000c)
`define MBOX_CSR_MBOX_DLEN                                                                          (32'hc)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_DATAIN                                                       (32'h30020010)
`define MBOX_CSR_MBOX_DATAIN                                                                        (32'h10)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_DATAOUT                                                      (32'h30020014)
`define MBOX_CSR_MBOX_DATAOUT                                                                       (32'h14)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_EXECUTE                                                      (32'h30020018)
`define MBOX_CSR_MBOX_EXECUTE                                                                       (32'h18)
`define MBOX_CSR_MBOX_EXECUTE_EXECUTE_LOW                                                           (0)
`define MBOX_CSR_MBOX_EXECUTE_EXECUTE_MASK                                                          (32'h1)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_STATUS                                                       (32'h3002001c)
`define MBOX_CSR_MBOX_STATUS                                                                        (32'h1c)
`define MBOX_CSR_MBOX_STATUS_STATUS_LOW                                                             (0)
`define MBOX_CSR_MBOX_STATUS_STATUS_MASK                                                            (32'hf)
`define MBOX_CSR_MBOX_STATUS_ECC_SINGLE_ERROR_LOW                                                   (4)
`define MBOX_CSR_MBOX_STATUS_ECC_SINGLE_ERROR_MASK                                                  (32'h10)
`define MBOX_CSR_MBOX_STATUS_ECC_DOUBLE_ERROR_LOW                                                   (5)
`define MBOX_CSR_MBOX_STATUS_ECC_DOUBLE_ERROR_MASK                                                  (32'h20)
`define MBOX_CSR_MBOX_STATUS_MBOX_FSM_PS_LOW                                                        (6)
`define MBOX_CSR_MBOX_STATUS_MBOX_FSM_PS_MASK                                                       (32'h1c0)
`define MBOX_CSR_MBOX_STATUS_SOC_HAS_LOCK_LOW                                                       (9)
`define MBOX_CSR_MBOX_STATUS_SOC_HAS_LOCK_MASK                                                      (32'h200)
`define MBOX_CSR_MBOX_STATUS_MBOX_RDPTR_LOW                                                         (10)
`define MBOX_CSR_MBOX_STATUS_MBOX_RDPTR_MASK                                                        (32'h1fffc00)
`define CALIPTRA_TOP_REG_MBOX_CSR_MBOX_UNLOCK                                                       (32'h30020020)
`define MBOX_CSR_MBOX_UNLOCK                                                                        (32'h20)
`define MBOX_CSR_MBOX_UNLOCK_UNLOCK_LOW                                                             (0)
`define MBOX_CSR_MBOX_UNLOCK_UNLOCK_MASK                                                            (32'h1)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_BASE_ADDR                                                   (32'h30021000)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_LOCK                                                        (32'h30021000)
`define SHA512_ACC_CSR_LOCK                                                                         (32'h0)
`define SHA512_ACC_CSR_LOCK_LOCK_LOW                                                                (0)
`define SHA512_ACC_CSR_LOCK_LOCK_MASK                                                               (32'h1)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_USER                                                        (32'h30021004)
`define SHA512_ACC_CSR_USER                                                                         (32'h4)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_MODE                                                        (32'h30021008)
`define SHA512_ACC_CSR_MODE                                                                         (32'h8)
`define SHA512_ACC_CSR_MODE_MODE_LOW                                                                (0)
`define SHA512_ACC_CSR_MODE_MODE_MASK                                                               (32'h3)
`define SHA512_ACC_CSR_MODE_ENDIAN_TOGGLE_LOW                                                       (2)
`define SHA512_ACC_CSR_MODE_ENDIAN_TOGGLE_MASK                                                      (32'h4)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_START_ADDRESS                                               (32'h3002100c)
`define SHA512_ACC_CSR_START_ADDRESS                                                                (32'hc)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DLEN                                                        (32'h30021010)
`define SHA512_ACC_CSR_DLEN                                                                         (32'h10)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DATAIN                                                      (32'h30021014)
`define SHA512_ACC_CSR_DATAIN                                                                       (32'h14)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_EXECUTE                                                     (32'h30021018)
`define SHA512_ACC_CSR_EXECUTE                                                                      (32'h18)
`define SHA512_ACC_CSR_EXECUTE_EXECUTE_LOW                                                          (0)
`define SHA512_ACC_CSR_EXECUTE_EXECUTE_MASK                                                         (32'h1)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_STATUS                                                      (32'h3002101c)
`define SHA512_ACC_CSR_STATUS                                                                       (32'h1c)
`define SHA512_ACC_CSR_STATUS_VALID_LOW                                                             (0)
`define SHA512_ACC_CSR_STATUS_VALID_MASK                                                            (32'h1)
`define SHA512_ACC_CSR_STATUS_SOC_HAS_LOCK_LOW                                                      (1)
`define SHA512_ACC_CSR_STATUS_SOC_HAS_LOCK_MASK                                                     (32'h2)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_0                                                    (32'h30021020)
`define SHA512_ACC_CSR_DIGEST_0                                                                     (32'h20)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_1                                                    (32'h30021024)
`define SHA512_ACC_CSR_DIGEST_1                                                                     (32'h24)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_2                                                    (32'h30021028)
`define SHA512_ACC_CSR_DIGEST_2                                                                     (32'h28)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_3                                                    (32'h3002102c)
`define SHA512_ACC_CSR_DIGEST_3                                                                     (32'h2c)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_4                                                    (32'h30021030)
`define SHA512_ACC_CSR_DIGEST_4                                                                     (32'h30)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_5                                                    (32'h30021034)
`define SHA512_ACC_CSR_DIGEST_5                                                                     (32'h34)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_6                                                    (32'h30021038)
`define SHA512_ACC_CSR_DIGEST_6                                                                     (32'h38)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_7                                                    (32'h3002103c)
`define SHA512_ACC_CSR_DIGEST_7                                                                     (32'h3c)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_8                                                    (32'h30021040)
`define SHA512_ACC_CSR_DIGEST_8                                                                     (32'h40)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_9                                                    (32'h30021044)
`define SHA512_ACC_CSR_DIGEST_9                                                                     (32'h44)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_10                                                   (32'h30021048)
`define SHA512_ACC_CSR_DIGEST_10                                                                    (32'h48)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_11                                                   (32'h3002104c)
`define SHA512_ACC_CSR_DIGEST_11                                                                    (32'h4c)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_12                                                   (32'h30021050)
`define SHA512_ACC_CSR_DIGEST_12                                                                    (32'h50)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_13                                                   (32'h30021054)
`define SHA512_ACC_CSR_DIGEST_13                                                                    (32'h54)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_14                                                   (32'h30021058)
`define SHA512_ACC_CSR_DIGEST_14                                                                    (32'h58)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_DIGEST_15                                                   (32'h3002105c)
`define SHA512_ACC_CSR_DIGEST_15                                                                    (32'h5c)
`define CALIPTRA_TOP_REG_SHA512_ACC_CSR_CONTROL                                                     (32'h30021060)
`define SHA512_ACC_CSR_CONTROL                                                                      (32'h60)
`define SHA512_ACC_CSR_CONTROL_ZEROIZE_LOW                                                          (0)
`define SHA512_ACC_CSR_CONTROL_ZEROIZE_MASK                                                         (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_BASE_ADDR                                             (32'h30030000)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL                                  (32'h30030000)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL                                                   (32'h0)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL_ICCM_ECC_UNC_LOW                                  (0)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL_ICCM_ECC_UNC_MASK                                 (32'h1)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL_DCCM_ECC_UNC_LOW                                  (1)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL_DCCM_ECC_UNC_MASK                                 (32'h2)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL_NMI_PIN_LOW                                       (2)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_FATAL_NMI_PIN_MASK                                      (32'h4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL                              (32'h30030004)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL                                               (32'h4)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_PROT_NO_LOCK_LOW                         (0)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_PROT_NO_LOCK_MASK                        (32'h1)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_PROT_OOO_LOW                             (1)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_PROT_OOO_MASK                            (32'h2)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_ECC_UNC_LOW                              (2)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_NON_FATAL_MBOX_ECC_UNC_MASK                             (32'h4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_FATAL                                  (32'h30030008)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_FATAL                                                   (32'h8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_NON_FATAL                              (32'h3003000c)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_NON_FATAL                                               (32'hc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_ENC                                    (32'h30030010)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_ERROR_ENC                                                     (32'h10)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_ENC                                    (32'h30030014)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_ERROR_ENC                                                     (32'h14)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                        (32'h30030018)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                         (32'h18)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                        (32'h3003001c)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                         (32'h1c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                        (32'h30030020)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                         (32'h20)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                        (32'h30030024)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                         (32'h24)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                        (32'h30030028)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                         (32'h28)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                        (32'h3003002c)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                         (32'h2c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                        (32'h30030030)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                         (32'h30)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                        (32'h30030034)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                         (32'h34)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_BOOT_STATUS                                     (32'h30030038)
`define GENERIC_AND_FUSE_REG_CPTRA_BOOT_STATUS                                                      (32'h38)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS                                     (32'h3003003c)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS                                                      (32'h3c)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_STATUS_LOW                                           (0)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_STATUS_MASK                                          (32'hffffff)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_IDEVID_CSR_READY_LOW                                 (24)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_IDEVID_CSR_READY_MASK                                (32'h1000000)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_BOOT_FSM_PS_LOW                                      (25)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_BOOT_FSM_PS_MASK                                     (32'he000000)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_READY_FOR_FW_LOW                                     (28)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_READY_FOR_FW_MASK                                    (32'h10000000)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_READY_FOR_RUNTIME_LOW                                (29)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_READY_FOR_RUNTIME_MASK                               (32'h20000000)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_READY_FOR_FUSES_LOW                                  (30)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_READY_FOR_FUSES_MASK                                 (32'h40000000)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_MAILBOX_FLOW_DONE_LOW                                (31)
`define GENERIC_AND_FUSE_REG_CPTRA_FLOW_STATUS_MAILBOX_FLOW_DONE_MASK                               (32'h80000000)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_RESET_REASON                                    (32'h30030040)
`define GENERIC_AND_FUSE_REG_CPTRA_RESET_REASON                                                     (32'h40)
`define GENERIC_AND_FUSE_REG_CPTRA_RESET_REASON_FW_UPD_RESET_LOW                                    (0)
`define GENERIC_AND_FUSE_REG_CPTRA_RESET_REASON_FW_UPD_RESET_MASK                                   (32'h1)
`define GENERIC_AND_FUSE_REG_CPTRA_RESET_REASON_WARM_RESET_LOW                                      (1)
`define GENERIC_AND_FUSE_REG_CPTRA_RESET_REASON_WARM_RESET_MASK                                     (32'h2)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE                                  (32'h30030044)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE                                                   (32'h44)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE_DEVICE_LIFECYCLE_LOW                              (0)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE_DEVICE_LIFECYCLE_MASK                             (32'h3)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE_DEBUG_LOCKED_LOW                                  (2)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE_DEBUG_LOCKED_MASK                                 (32'h4)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE_SCAN_MODE_LOW                                     (3)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE_SCAN_MODE_MASK                                    (32'h8)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE_RSVD_LOW                                          (4)
`define GENERIC_AND_FUSE_REG_CPTRA_SECURITY_STATE_RSVD_MASK                                         (32'hfffffff0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_0                             (32'h30030048)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_0                                              (32'h48)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_1                             (32'h3003004c)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_1                                              (32'h4c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_2                             (32'h30030050)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_2                                              (32'h50)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_3                             (32'h30030054)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_3                                              (32'h54)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_4                             (32'h30030058)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_VALID_PAUSER_4                                              (32'h58)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_0                              (32'h3003005c)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_0                                               (32'h5c)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_0_LOCK_LOW                                      (0)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_0_LOCK_MASK                                     (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_1                              (32'h30030060)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_1                                               (32'h60)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_1_LOCK_LOW                                      (0)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_1_LOCK_MASK                                     (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_2                              (32'h30030064)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_2                                               (32'h64)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_2_LOCK_LOW                                      (0)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_2_LOCK_MASK                                     (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_3                              (32'h30030068)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_3                                               (32'h68)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_3_LOCK_LOW                                      (0)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_3_LOCK_MASK                                     (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_4                              (32'h3003006c)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_4                                               (32'h6c)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_4_LOCK_LOW                                      (0)
`define GENERIC_AND_FUSE_REG_CPTRA_MBOX_PAUSER_LOCK_4_LOCK_MASK                                     (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_VALID_PAUSER                               (32'h30030070)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_VALID_PAUSER                                                (32'h70)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_PAUSER_LOCK                                (32'h30030074)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_PAUSER_LOCK                                                 (32'h74)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_PAUSER_LOCK_LOCK_LOW                                        (0)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_PAUSER_LOCK_LOCK_MASK                                       (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_0                                     (32'h30030078)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_0                                                      (32'h78)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_1                                     (32'h3003007c)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_1                                                      (32'h7c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_2                                     (32'h30030080)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_2                                                      (32'h80)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_3                                     (32'h30030084)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_3                                                      (32'h84)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_4                                     (32'h30030088)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_4                                                      (32'h88)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_5                                     (32'h3003008c)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_5                                                      (32'h8c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_6                                     (32'h30030090)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_6                                                      (32'h90)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_7                                     (32'h30030094)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_7                                                      (32'h94)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_8                                     (32'h30030098)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_8                                                      (32'h98)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_9                                     (32'h3003009c)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_9                                                      (32'h9c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_10                                    (32'h300300a0)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_10                                                     (32'ha0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_11                                    (32'h300300a4)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_DATA_11                                                     (32'ha4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_CTRL                                       (32'h300300a8)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_CTRL                                                        (32'ha8)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_CTRL_CLEAR_LOW                                              (0)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_CTRL_CLEAR_MASK                                             (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TRNG_STATUS                                     (32'h300300ac)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_STATUS                                                      (32'hac)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_STATUS_DATA_REQ_LOW                                         (0)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_STATUS_DATA_REQ_MASK                                        (32'h1)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_STATUS_DATA_WR_DONE_LOW                                     (1)
`define GENERIC_AND_FUSE_REG_CPTRA_TRNG_STATUS_DATA_WR_DONE_MASK                                    (32'h2)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FUSE_WR_DONE                                    (32'h300300b0)
`define GENERIC_AND_FUSE_REG_CPTRA_FUSE_WR_DONE                                                     (32'hb0)
`define GENERIC_AND_FUSE_REG_CPTRA_FUSE_WR_DONE_DONE_LOW                                            (0)
`define GENERIC_AND_FUSE_REG_CPTRA_FUSE_WR_DONE_DONE_MASK                                           (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_TIMER_CONFIG                                    (32'h300300b4)
`define GENERIC_AND_FUSE_REG_CPTRA_TIMER_CONFIG                                                     (32'hb4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_BOOTFSM_GO                                      (32'h300300b8)
`define GENERIC_AND_FUSE_REG_CPTRA_BOOTFSM_GO                                                       (32'hb8)
`define GENERIC_AND_FUSE_REG_CPTRA_BOOTFSM_GO_GO_LOW                                                (0)
`define GENERIC_AND_FUSE_REG_CPTRA_BOOTFSM_GO_GO_MASK                                               (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_DBG_MANUF_SERVICE_REG                           (32'h300300bc)
`define GENERIC_AND_FUSE_REG_CPTRA_DBG_MANUF_SERVICE_REG                                            (32'hbc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_CLK_GATING_EN                                   (32'h300300c0)
`define GENERIC_AND_FUSE_REG_CPTRA_CLK_GATING_EN                                                    (32'hc0)
`define GENERIC_AND_FUSE_REG_CPTRA_CLK_GATING_EN_CLK_GATING_EN_LOW                                  (0)
`define GENERIC_AND_FUSE_REG_CPTRA_CLK_GATING_EN_CLK_GATING_EN_MASK                                 (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_GENERIC_INPUT_WIRES_0                           (32'h300300c4)
`define GENERIC_AND_FUSE_REG_CPTRA_GENERIC_INPUT_WIRES_0                                            (32'hc4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_GENERIC_INPUT_WIRES_1                           (32'h300300c8)
`define GENERIC_AND_FUSE_REG_CPTRA_GENERIC_INPUT_WIRES_1                                            (32'hc8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                          (32'h300300cc)
`define GENERIC_AND_FUSE_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                           (32'hcc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                          (32'h300300d0)
`define GENERIC_AND_FUSE_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                           (32'hd0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_REV_ID                                       (32'h300300d4)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_REV_ID                                                        (32'hd4)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_REV_ID_CPTRA_GENERATION_LOW                                   (0)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_REV_ID_CPTRA_GENERATION_MASK                                  (32'hffff)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_REV_ID_SOC_STEPPING_ID_LOW                                    (16)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_REV_ID_SOC_STEPPING_ID_MASK                                   (32'hffff0000)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_REV_ID_0                                     (32'h300300d8)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_REV_ID_0                                                      (32'hd8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FW_REV_ID_1                                     (32'h300300dc)
`define GENERIC_AND_FUSE_REG_CPTRA_FW_REV_ID_1                                                      (32'hdc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG                                       (32'h300300e0)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG                                                        (32'he0)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_ITRNG_EN_LOW                                           (0)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_ITRNG_EN_MASK                                          (32'h1)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_QSPI_EN_LOW                                            (1)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_QSPI_EN_MASK                                           (32'h2)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_I3C_EN_LOW                                             (2)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_I3C_EN_MASK                                            (32'h4)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_UART_EN_LOW                                            (3)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_UART_EN_MASK                                           (32'h8)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_LMS_ACC_EN_LOW                                         (4)
`define GENERIC_AND_FUSE_REG_CPTRA_HW_CONFIG_LMS_ACC_EN_MASK                                        (32'h10)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_EN                                   (32'h300300e4)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_EN                                                    (32'he4)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_EN_TIMER1_EN_LOW                                      (0)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_EN_TIMER1_EN_MASK                                     (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_CTRL                                 (32'h300300e8)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_CTRL                                                  (32'he8)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_CTRL_TIMER1_RESTART_LOW                               (0)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_CTRL_TIMER1_RESTART_MASK                              (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_0                     (32'h300300ec)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_0                                      (32'hec)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_1                     (32'h300300f0)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_1                                      (32'hf0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_EN                                   (32'h300300f4)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_EN                                                    (32'hf4)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_EN_TIMER2_EN_LOW                                      (0)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_EN_TIMER2_EN_MASK                                     (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_CTRL                                 (32'h300300f8)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_CTRL                                                  (32'hf8)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_CTRL_TIMER2_RESTART_LOW                               (0)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_CTRL_TIMER2_RESTART_MASK                              (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_0                     (32'h300300fc)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_0                                      (32'hfc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_1                     (32'h30030100)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_1                                      (32'h100)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_STATUS                                      (32'h30030104)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_STATUS                                                       (32'h104)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_STATUS_T1_TIMEOUT_LOW                                        (0)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_STATUS_T1_TIMEOUT_MASK                                       (32'h1)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_STATUS_T2_TIMEOUT_LOW                                        (1)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_STATUS_T2_TIMEOUT_MASK                                       (32'h2)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FUSE_VALID_PAUSER                               (32'h30030108)
`define GENERIC_AND_FUSE_REG_CPTRA_FUSE_VALID_PAUSER                                                (32'h108)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_FUSE_PAUSER_LOCK                                (32'h3003010c)
`define GENERIC_AND_FUSE_REG_CPTRA_FUSE_PAUSER_LOCK                                                 (32'h10c)
`define GENERIC_AND_FUSE_REG_CPTRA_FUSE_PAUSER_LOCK_LOCK_LOW                                        (0)
`define GENERIC_AND_FUSE_REG_CPTRA_FUSE_PAUSER_LOCK_LOCK_MASK                                       (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_CFG_0                                       (32'h30030110)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_CFG_0                                                        (32'h110)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_WDT_CFG_1                                       (32'h30030114)
`define GENERIC_AND_FUSE_REG_CPTRA_WDT_CFG_1                                                        (32'h114)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0                          (32'h30030118)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0                                           (32'h118)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0_LOW_THRESHOLD_LOW                         (0)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0_LOW_THRESHOLD_MASK                        (32'hffff)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0_HIGH_THRESHOLD_LOW                        (16)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0_HIGH_THRESHOLD_MASK                       (32'hffff0000)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1                          (32'h3003011c)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1                                           (32'h11c)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1_REPETITION_COUNT_LOW                      (0)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1_REPETITION_COUNT_MASK                     (32'hffff)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1_RSVD_LOW                                  (16)
`define GENERIC_AND_FUSE_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1_RSVD_MASK                                 (32'hffff0000)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_RSVD_REG_0                                      (32'h30030120)
`define GENERIC_AND_FUSE_REG_CPTRA_RSVD_REG_0                                                       (32'h120)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_CPTRA_RSVD_REG_1                                      (32'h30030124)
`define GENERIC_AND_FUSE_REG_CPTRA_RSVD_REG_1                                                       (32'h124)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_0                                       (32'h30030200)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_0                                                        (32'h200)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_1                                       (32'h30030204)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_1                                                        (32'h204)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_2                                       (32'h30030208)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_2                                                        (32'h208)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_3                                       (32'h3003020c)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_3                                                        (32'h20c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_4                                       (32'h30030210)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_4                                                        (32'h210)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_5                                       (32'h30030214)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_5                                                        (32'h214)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_6                                       (32'h30030218)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_6                                                        (32'h218)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_7                                       (32'h3003021c)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_7                                                        (32'h21c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_8                                       (32'h30030220)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_8                                                        (32'h220)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_9                                       (32'h30030224)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_9                                                        (32'h224)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_10                                      (32'h30030228)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_10                                                       (32'h228)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_11                                      (32'h3003022c)
`define GENERIC_AND_FUSE_REG_FUSE_UDS_SEED_11                                                       (32'h22c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_0                                  (32'h30030230)
`define GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_0                                                   (32'h230)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_1                                  (32'h30030234)
`define GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_1                                                   (32'h234)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_2                                  (32'h30030238)
`define GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_2                                                   (32'h238)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_3                                  (32'h3003023c)
`define GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_3                                                   (32'h23c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_4                                  (32'h30030240)
`define GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_4                                                   (32'h240)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_5                                  (32'h30030244)
`define GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_5                                                   (32'h244)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_6                                  (32'h30030248)
`define GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_6                                                   (32'h248)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_7                                  (32'h3003024c)
`define GENERIC_AND_FUSE_REG_FUSE_FIELD_ENTROPY_7                                                   (32'h24c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_0                           (32'h30030250)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_0                                            (32'h250)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_1                           (32'h30030254)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_1                                            (32'h254)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_2                           (32'h30030258)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_2                                            (32'h258)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_3                           (32'h3003025c)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_3                                            (32'h25c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_4                           (32'h30030260)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_4                                            (32'h260)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_5                           (32'h30030264)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_5                                            (32'h264)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_6                           (32'h30030268)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_6                                            (32'h268)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_7                           (32'h3003026c)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_7                                            (32'h26c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_8                           (32'h30030270)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_8                                            (32'h270)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_9                           (32'h30030274)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_9                                            (32'h274)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_10                          (32'h30030278)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_10                                           (32'h278)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_11                          (32'h3003027c)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_11                                           (32'h27c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK                        (32'h30030280)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK                                         (32'h280)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK_MASK_LOW                                (0)
`define GENERIC_AND_FUSE_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK_MASK_MASK                               (32'hf)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_0                                  (32'h30030284)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_0                                                   (32'h284)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_1                                  (32'h30030288)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_1                                                   (32'h288)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_2                                  (32'h3003028c)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_2                                                   (32'h28c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_3                                  (32'h30030290)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_3                                                   (32'h290)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_4                                  (32'h30030294)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_4                                                   (32'h294)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_5                                  (32'h30030298)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_5                                                   (32'h298)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_6                                  (32'h3003029c)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_6                                                   (32'h29c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_7                                  (32'h300302a0)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_7                                                   (32'h2a0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_8                                  (32'h300302a4)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_8                                                   (32'h2a4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_9                                  (32'h300302a8)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_9                                                   (32'h2a8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_10                                 (32'h300302ac)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_10                                                  (32'h2ac)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_11                                 (32'h300302b0)
`define GENERIC_AND_FUSE_REG_FUSE_OWNER_PK_HASH_11                                                  (32'h2b0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_FMC_KEY_MANIFEST_SVN                             (32'h300302b4)
`define GENERIC_AND_FUSE_REG_FUSE_FMC_KEY_MANIFEST_SVN                                              (32'h2b4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_0                                    (32'h300302b8)
`define GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_0                                                     (32'h2b8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_1                                    (32'h300302bc)
`define GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_1                                                     (32'h2bc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_2                                    (32'h300302c0)
`define GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_2                                                     (32'h2c0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_3                                    (32'h300302c4)
`define GENERIC_AND_FUSE_REG_FUSE_RUNTIME_SVN_3                                                     (32'h2c4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_ANTI_ROLLBACK_DISABLE                            (32'h300302c8)
`define GENERIC_AND_FUSE_REG_FUSE_ANTI_ROLLBACK_DISABLE                                             (32'h2c8)
`define GENERIC_AND_FUSE_REG_FUSE_ANTI_ROLLBACK_DISABLE_DIS_LOW                                     (0)
`define GENERIC_AND_FUSE_REG_FUSE_ANTI_ROLLBACK_DISABLE_DIS_MASK                                    (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_0                               (32'h300302cc)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_0                                                (32'h2cc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_1                               (32'h300302d0)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_1                                                (32'h2d0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_2                               (32'h300302d4)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_2                                                (32'h2d4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_3                               (32'h300302d8)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_3                                                (32'h2d8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_4                               (32'h300302dc)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_4                                                (32'h2dc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_5                               (32'h300302e0)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_5                                                (32'h2e0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_6                               (32'h300302e4)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_6                                                (32'h2e4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_7                               (32'h300302e8)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_7                                                (32'h2e8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_8                               (32'h300302ec)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_8                                                (32'h2ec)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_9                               (32'h300302f0)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_9                                                (32'h2f0)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_10                              (32'h300302f4)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_10                                               (32'h2f4)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_11                              (32'h300302f8)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_11                                               (32'h2f8)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_12                              (32'h300302fc)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_12                                               (32'h2fc)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_13                              (32'h30030300)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_13                                               (32'h300)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_14                              (32'h30030304)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_14                                               (32'h304)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_15                              (32'h30030308)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_15                                               (32'h308)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_16                              (32'h3003030c)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_16                                               (32'h30c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_17                              (32'h30030310)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_17                                               (32'h310)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_18                              (32'h30030314)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_18                                               (32'h314)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_19                              (32'h30030318)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_19                                               (32'h318)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_20                              (32'h3003031c)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_20                                               (32'h31c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_21                              (32'h30030320)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_21                                               (32'h320)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_22                              (32'h30030324)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_22                                               (32'h324)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_23                              (32'h30030328)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_CERT_ATTR_23                                               (32'h328)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_0                            (32'h3003032c)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                             (32'h32c)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_1                            (32'h30030330)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                             (32'h330)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_2                            (32'h30030334)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                             (32'h334)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_3                            (32'h30030338)
`define GENERIC_AND_FUSE_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                             (32'h338)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_LIFE_CYCLE                                       (32'h3003033c)
`define GENERIC_AND_FUSE_REG_FUSE_LIFE_CYCLE                                                        (32'h33c)
`define GENERIC_AND_FUSE_REG_FUSE_LIFE_CYCLE_LIFE_CYCLE_LOW                                         (0)
`define GENERIC_AND_FUSE_REG_FUSE_LIFE_CYCLE_LIFE_CYCLE_MASK                                        (32'h3)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_LMS_VERIFY                                       (32'h30030340)
`define GENERIC_AND_FUSE_REG_FUSE_LMS_VERIFY                                                        (32'h340)
`define GENERIC_AND_FUSE_REG_FUSE_LMS_VERIFY_LMS_VERIFY_LOW                                         (0)
`define GENERIC_AND_FUSE_REG_FUSE_LMS_VERIFY_LMS_VERIFY_MASK                                        (32'h1)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_LMS_REVOCATION                                   (32'h30030344)
`define GENERIC_AND_FUSE_REG_FUSE_LMS_REVOCATION                                                    (32'h344)
`define CALIPTRA_TOP_REG_GENERIC_AND_FUSE_REG_FUSE_SOC_STEPPING_ID                                  (32'h30030348)
`define GENERIC_AND_FUSE_REG_FUSE_SOC_STEPPING_ID                                                   (32'h348)
`define GENERIC_AND_FUSE_REG_FUSE_SOC_STEPPING_ID_SOC_STEPPING_ID_LOW                               (0)
`define GENERIC_AND_FUSE_REG_FUSE_SOC_STEPPING_ID_SOC_STEPPING_ID_MASK                              (32'hffff)


`endif