// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Write enable and data arbitration logic for register slice conforming to Comportibility guide.

module caliptra_prim_subreg_arb
  import caliptra_prim_subreg_pkg::*;
#(
  parameter int         DW       = 32,
  parameter sw_access_e SwAccess = SwAccessRW,
  parameter bit         Mubi     = 1'b0
) (
  // From SW: valid for RW, WO, W1C, W1S, W0C, RC.
  // In case of RC, top connects read pulse to we.
  input          we,
  input [DW-1:0] wd,

  // From HW: valid for HRW, HWO.
  input          de,
  input [DW-1:0] d,

  // From register: actual reg value.
  input [DW-1:0] q,

  // To register: actual write enable and write data.
  output logic          wr_en,
  output logic [DW-1:0] wr_data
);
  import caliptra_prim_mubi_pkg::*;
  import caliptra_prim_mubi_pkg::*;

  if (SwAccess inside {SwAccessRW, SwAccessWO}) begin : gen_w
    assign wr_en   = we | de;
    assign wr_data = (we == 1'b1) ? wd : d; // SW higher priority
    // Unused q - Prevent lint errors.
    logic [DW-1:0] unused_q;
    //VCS coverage off
    // pragma coverage off
    //VCS coverage off
    // pragma coverage off
    assign unused_q = q;
    //VCS coverage on
    // pragma coverage on
    //VCS coverage on
    // pragma coverage on
  end else if (SwAccess == SwAccessRO) begin : gen_ro
    assign wr_en   = de;
    assign wr_data = d;
    // Unused we, wd, q - Prevent lint errors.
    logic          unused_we;
    logic [DW-1:0] unused_wd;
    logic [DW-1:0] unused_q;
    //VCS coverage off
    // pragma coverage off
    //VCS coverage off
    // pragma coverage off
    assign unused_we = we;
    assign unused_wd = wd;
    assign unused_q  = q;
    //VCS coverage on
    // pragma coverage on
    //VCS coverage on
    // pragma coverage on
  end else if (SwAccess == SwAccessW1S) begin : gen_w1s
    // If SwAccess is W1S, then assume hw tries to clear.
    // So, give a chance HW to clear when SW tries to set.
    // If both try to set/clr at the same bit pos, SW wins.
    assign wr_en   = we | de;
    if (Mubi) begin : gen_mubi
      if (DW == 4) begin : gen_mubi4
        assign wr_data = caliptra_prim_mubi_pkg::mubi4_or_hi(caliptra_prim_mubi_pkg::mubi4_t'(de ? d : q),
                                                             (we ? caliptra_prim_mubi_pkg::mubi4_t'(wd) :
                                                                   caliptra_prim_mubi_pkg::MuBi4False));
      end else if (DW == 8) begin : gen_mubi8
        assign wr_data = caliptra_prim_mubi_pkg::mubi8_or_hi(caliptra_prim_mubi_pkg::mubi8_t'(de ? d : q),
                                                             (we ? caliptra_prim_mubi_pkg::mubi8_t'(wd) :
                                                                   caliptra_prim_mubi_pkg::MuBi8False));
      end else if (DW == 12) begin : gen_mubi12
        assign wr_data = caliptra_prim_mubi_pkg::mubi12_or_hi(caliptra_prim_mubi_pkg::mubi12_t'(de ? d : q),
                                                              (we ? caliptra_prim_mubi_pkg::mubi12_t'(wd) :
                                                                    caliptra_prim_mubi_pkg::MuBi12False));
      end else if (DW == 16) begin : gen_mubi16
        assign wr_data = caliptra_prim_mubi_pkg::mubi16_or_hi(caliptra_prim_mubi_pkg::mubi16_t'(de ? d : q),
                                                              (we ? caliptra_prim_mubi_pkg::mubi16_t'(wd) :
                                                                    caliptra_prim_mubi_pkg::MuBi16False));
      end else begin : gen_invalid_mubi
        $error("%m: Invalid width for MuBi");
      end
    end else begin : gen_non_mubi
      assign wr_data = (de ? d : q) | (we ? wd : '0);
    end
  end else if (SwAccess == SwAccessW1C) begin : gen_w1c
    // If SwAccess is W1C, then assume hw tries to set.
    // So, give a chance HW to set when SW tries to clear.
    // If both try to set/clr at the same bit pos, SW wins.
    assign wr_en   = we | de;
    if (Mubi) begin : gen_mubi
      if (DW == 4) begin : gen_mubi4
        assign wr_data = caliptra_prim_mubi_pkg::mubi4_and_hi(caliptra_prim_mubi_pkg::mubi4_t'(de ? d : q),
                                                              (we ? caliptra_prim_mubi_pkg::mubi4_t'(~wd) :
                                                                    caliptra_prim_mubi_pkg::MuBi4True));
      end else if (DW == 8) begin : gen_mubi8
        assign wr_data = caliptra_prim_mubi_pkg::mubi8_and_hi(caliptra_prim_mubi_pkg::mubi8_t'(de ? d : q),
                                                              (we ? caliptra_prim_mubi_pkg::mubi8_t'(~wd) :
                                                                    caliptra_prim_mubi_pkg::MuBi8True));
      end else if (DW == 12) begin : gen_mubi12
        assign wr_data = caliptra_prim_mubi_pkg::mubi12_and_hi(caliptra_prim_mubi_pkg::mubi12_t'(de ? d : q),
                                                               (we ? caliptra_prim_mubi_pkg::mubi12_t'(~wd) :
                                                                     caliptra_prim_mubi_pkg::MuBi12True));
      end else if (DW == 16) begin : gen_mubi16
        assign wr_data = caliptra_prim_mubi_pkg::mubi16_and_hi(caliptra_prim_mubi_pkg::mubi16_t'(de ? d : q),
                                                               (we ? caliptra_prim_mubi_pkg::mubi16_t'(~wd) :
                                                                     caliptra_prim_mubi_pkg::MuBi16True));
      end else begin : gen_invalid_mubi
        $error("%m: Invalid width for MuBi");
      end
    end else begin : gen_non_mubi
      assign wr_data = (de ? d : q) & (we ? ~wd : '1);
    end
  end else if (SwAccess == SwAccessW0C) begin : gen_w0c
    assign wr_en   = we | de;
    if (Mubi) begin : gen_mubi
      if (DW == 4) begin : gen_mubi4
        assign wr_data = caliptra_prim_mubi_pkg::mubi4_and_hi(caliptra_prim_mubi_pkg::mubi4_t'(de ? d : q),
                                                              (we ? caliptra_prim_mubi_pkg::mubi4_t'(wd) :
                                                                    caliptra_prim_mubi_pkg::MuBi4True));
      end else if (DW == 8) begin : gen_mubi8
        assign wr_data = caliptra_prim_mubi_pkg::mubi8_and_hi(caliptra_prim_mubi_pkg::mubi8_t'(de ? d : q),
                                                              (we ? caliptra_prim_mubi_pkg::mubi8_t'(wd) :
                                                                    caliptra_prim_mubi_pkg::MuBi8True));
      end else if (DW == 12) begin : gen_mubi12
        assign wr_data = caliptra_prim_mubi_pkg::mubi12_and_hi(caliptra_prim_mubi_pkg::mubi12_t'(de ? d : q),
                                                               (we ? caliptra_prim_mubi_pkg::mubi12_t'(wd) :
                                                                     caliptra_prim_mubi_pkg::MuBi12True));
      end else if (DW == 16) begin : gen_mubi16
        assign wr_data = caliptra_prim_mubi_pkg::mubi16_and_hi(caliptra_prim_mubi_pkg::mubi16_t'(de ? d : q),
                                                               (we ? caliptra_prim_mubi_pkg::mubi16_t'(wd) :
                                                                     caliptra_prim_mubi_pkg::MuBi16True));
      end else begin : gen_invalid_mubi
        $error("%m: Invalid width for MuBi");
      end
    end else begin : gen_non_mubi
      assign wr_data = (de ? d : q) & (we ? wd : '1);
    end
  end else if (SwAccess == SwAccessRC) begin : gen_rc
    // This swtype is not recommended but exists for compatibility.
    // WARN: we signal is actually read signal not write enable.
    assign wr_en  = we | de;
    if (Mubi) begin : gen_mubi
      if (DW == 4) begin : gen_mubi4
        assign wr_data = caliptra_prim_mubi_pkg::mubi4_and_hi(caliptra_prim_mubi_pkg::mubi4_t'(de ? d : q),
                                                              (we ? caliptra_prim_mubi_pkg::MuBi4False :
                                                                    caliptra_prim_mubi_pkg::MuBi4True));
      end else if (DW == 8) begin : gen_mubi8
        assign wr_data = caliptra_prim_mubi_pkg::mubi8_and_hi(caliptra_prim_mubi_pkg::mubi8_t'(de ? d : q),
                                                              (we ? caliptra_prim_mubi_pkg::MuBi8False :
                                                                    caliptra_prim_mubi_pkg::MuBi8True));
      end else if (DW == 12) begin : gen_mubi12
        assign wr_data = caliptra_prim_mubi_pkg::mubi12_and_hi(caliptra_prim_mubi_pkg::mubi12_t'(de ? d : q),
                                                               (we ? caliptra_prim_mubi_pkg::MuBi12False :
                                                                     caliptra_prim_mubi_pkg::MuBi12True));
      end else if (DW == 16) begin : gen_mubi16
        assign wr_data = caliptra_prim_mubi_pkg::mubi16_and_hi(caliptra_prim_mubi_pkg::mubi16_t'(de ? d : q),
                                                               (we ? caliptra_prim_mubi_pkg::mubi16_t'(wd) :
                                                                     caliptra_prim_mubi_pkg::MuBi16True));
      end else begin : gen_invalid_mubi
        $error("%m: Invalid width for MuBi");
      end
    end else begin : gen_non_mubi
      assign wr_data = (de ? d : q) & (we ? '0 : '1);
    end
    // Unused wd - Prevent lint errors.
    logic [DW-1:0] unused_wd;
    //VCS coverage off
    // pragma coverage off
    //VCS coverage off
    // pragma coverage off
    assign unused_wd = wd;
    //VCS coverage on
    // pragma coverage on
    //VCS coverage on
    // pragma coverage on
  end else begin : gen_hw
    assign wr_en   = de;
    assign wr_data = d;
    // Unused we, wd, q - Prevent lint errors.
    logic          unused_we;
    logic [DW-1:0] unused_wd;
    logic [DW-1:0] unused_q;
    //VCS coverage off
    // pragma coverage off
    //VCS coverage off
    // pragma coverage off
    assign unused_we = we;
    assign unused_wd = wd;
    assign unused_q  = q;
    //VCS coverage on
    // pragma coverage on
    //VCS coverage on
    // pragma coverage on
  end

endmodule
