//
// File: hvl_qvip_ahb_lite_slave.sv
//
// Generated from Mentor VIP Configurator (20220406)
// Generated using Mentor VIP Library ( 2022.2 : 04/20/2022:16:06 )
//
module hvl_qvip_ahb_lite_slave;
    import uvm_pkg::*;
    
    `include "test_packages.svh"
    
    initial
    begin
        run_test();
    end

endmodule: hvl_qvip_ahb_lite_slave
