// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef CALIPTRA_REG_DEFINES_HEADER
`define CALIPTRA_REG_DEFINES_HEADER


`define CLP_BASE_ADDR                                                                               (32'h0)
`define CLP_DOE_REG_BASE_ADDR                                                                       (32'h10000000)
`define CLP_DOE_REG_DOE_IV_0                                                                        (32'h10000000)
`define CLP_DOE_REG_DOE_IV_1                                                                        (32'h10000004)
`define CLP_DOE_REG_DOE_IV_2                                                                        (32'h10000008)
`define CLP_DOE_REG_DOE_IV_3                                                                        (32'h1000000c)
`define CLP_DOE_REG_DOE_CTRL                                                                        (32'h10000010)
`define CLP_DOE_REG_DOE_STATUS                                                                      (32'h10000014)
`define CLP_DOE_REG_INTR_BLOCK_RF_START                                                             (32'h10000800)
`define CLP_DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10000800)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10000804)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10000808)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1000080c)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10000810)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10000814)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10000818)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1000081c)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10000820)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                               (32'h10000900)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                               (32'h10000904)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                               (32'h10000908)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                               (32'h1000090c)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10000980)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                          (32'h10000a00)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                          (32'h10000a04)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                          (32'h10000a08)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                          (32'h10000a0c)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10000a10)
`define CLP_ECC_REG_BASE_ADDR                                                                       (32'h10008000)
`define CLP_ECC_REG_ECC_NAME_0                                                                      (32'h10008000)
`define CLP_ECC_REG_ECC_NAME_1                                                                      (32'h10008004)
`define CLP_ECC_REG_ECC_VERSION_0                                                                   (32'h10008008)
`define CLP_ECC_REG_ECC_VERSION_1                                                                   (32'h1000800c)
`define CLP_ECC_REG_ECC_CTRL                                                                        (32'h10008010)
`define CLP_ECC_REG_ECC_STATUS                                                                      (32'h10008018)
`define CLP_ECC_REG_ECC_SEED_0                                                                      (32'h10008080)
`define CLP_ECC_REG_ECC_SEED_1                                                                      (32'h10008084)
`define CLP_ECC_REG_ECC_SEED_2                                                                      (32'h10008088)
`define CLP_ECC_REG_ECC_SEED_3                                                                      (32'h1000808c)
`define CLP_ECC_REG_ECC_SEED_4                                                                      (32'h10008090)
`define CLP_ECC_REG_ECC_SEED_5                                                                      (32'h10008094)
`define CLP_ECC_REG_ECC_SEED_6                                                                      (32'h10008098)
`define CLP_ECC_REG_ECC_SEED_7                                                                      (32'h1000809c)
`define CLP_ECC_REG_ECC_SEED_8                                                                      (32'h100080a0)
`define CLP_ECC_REG_ECC_SEED_9                                                                      (32'h100080a4)
`define CLP_ECC_REG_ECC_SEED_10                                                                     (32'h100080a8)
`define CLP_ECC_REG_ECC_SEED_11                                                                     (32'h100080ac)
`define CLP_ECC_REG_ECC_MSG_0                                                                       (32'h10008100)
`define CLP_ECC_REG_ECC_MSG_1                                                                       (32'h10008104)
`define CLP_ECC_REG_ECC_MSG_2                                                                       (32'h10008108)
`define CLP_ECC_REG_ECC_MSG_3                                                                       (32'h1000810c)
`define CLP_ECC_REG_ECC_MSG_4                                                                       (32'h10008110)
`define CLP_ECC_REG_ECC_MSG_5                                                                       (32'h10008114)
`define CLP_ECC_REG_ECC_MSG_6                                                                       (32'h10008118)
`define CLP_ECC_REG_ECC_MSG_7                                                                       (32'h1000811c)
`define CLP_ECC_REG_ECC_MSG_8                                                                       (32'h10008120)
`define CLP_ECC_REG_ECC_MSG_9                                                                       (32'h10008124)
`define CLP_ECC_REG_ECC_MSG_10                                                                      (32'h10008128)
`define CLP_ECC_REG_ECC_MSG_11                                                                      (32'h1000812c)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_0                                                               (32'h10008180)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_1                                                               (32'h10008184)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_2                                                               (32'h10008188)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_3                                                               (32'h1000818c)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_4                                                               (32'h10008190)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_5                                                               (32'h10008194)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_6                                                               (32'h10008198)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_7                                                               (32'h1000819c)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_8                                                               (32'h100081a0)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_9                                                               (32'h100081a4)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_10                                                              (32'h100081a8)
`define CLP_ECC_REG_ECC_PRIVKEY_OUT_11                                                              (32'h100081ac)
`define CLP_ECC_REG_ECC_PUBKEY_X_0                                                                  (32'h10008200)
`define CLP_ECC_REG_ECC_PUBKEY_X_1                                                                  (32'h10008204)
`define CLP_ECC_REG_ECC_PUBKEY_X_2                                                                  (32'h10008208)
`define CLP_ECC_REG_ECC_PUBKEY_X_3                                                                  (32'h1000820c)
`define CLP_ECC_REG_ECC_PUBKEY_X_4                                                                  (32'h10008210)
`define CLP_ECC_REG_ECC_PUBKEY_X_5                                                                  (32'h10008214)
`define CLP_ECC_REG_ECC_PUBKEY_X_6                                                                  (32'h10008218)
`define CLP_ECC_REG_ECC_PUBKEY_X_7                                                                  (32'h1000821c)
`define CLP_ECC_REG_ECC_PUBKEY_X_8                                                                  (32'h10008220)
`define CLP_ECC_REG_ECC_PUBKEY_X_9                                                                  (32'h10008224)
`define CLP_ECC_REG_ECC_PUBKEY_X_10                                                                 (32'h10008228)
`define CLP_ECC_REG_ECC_PUBKEY_X_11                                                                 (32'h1000822c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_0                                                                  (32'h10008280)
`define CLP_ECC_REG_ECC_PUBKEY_Y_1                                                                  (32'h10008284)
`define CLP_ECC_REG_ECC_PUBKEY_Y_2                                                                  (32'h10008288)
`define CLP_ECC_REG_ECC_PUBKEY_Y_3                                                                  (32'h1000828c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_4                                                                  (32'h10008290)
`define CLP_ECC_REG_ECC_PUBKEY_Y_5                                                                  (32'h10008294)
`define CLP_ECC_REG_ECC_PUBKEY_Y_6                                                                  (32'h10008298)
`define CLP_ECC_REG_ECC_PUBKEY_Y_7                                                                  (32'h1000829c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_8                                                                  (32'h100082a0)
`define CLP_ECC_REG_ECC_PUBKEY_Y_9                                                                  (32'h100082a4)
`define CLP_ECC_REG_ECC_PUBKEY_Y_10                                                                 (32'h100082a8)
`define CLP_ECC_REG_ECC_PUBKEY_Y_11                                                                 (32'h100082ac)
`define CLP_ECC_REG_ECC_SIGN_R_0                                                                    (32'h10008300)
`define CLP_ECC_REG_ECC_SIGN_R_1                                                                    (32'h10008304)
`define CLP_ECC_REG_ECC_SIGN_R_2                                                                    (32'h10008308)
`define CLP_ECC_REG_ECC_SIGN_R_3                                                                    (32'h1000830c)
`define CLP_ECC_REG_ECC_SIGN_R_4                                                                    (32'h10008310)
`define CLP_ECC_REG_ECC_SIGN_R_5                                                                    (32'h10008314)
`define CLP_ECC_REG_ECC_SIGN_R_6                                                                    (32'h10008318)
`define CLP_ECC_REG_ECC_SIGN_R_7                                                                    (32'h1000831c)
`define CLP_ECC_REG_ECC_SIGN_R_8                                                                    (32'h10008320)
`define CLP_ECC_REG_ECC_SIGN_R_9                                                                    (32'h10008324)
`define CLP_ECC_REG_ECC_SIGN_R_10                                                                   (32'h10008328)
`define CLP_ECC_REG_ECC_SIGN_R_11                                                                   (32'h1000832c)
`define CLP_ECC_REG_ECC_SIGN_S_0                                                                    (32'h10008380)
`define CLP_ECC_REG_ECC_SIGN_S_1                                                                    (32'h10008384)
`define CLP_ECC_REG_ECC_SIGN_S_2                                                                    (32'h10008388)
`define CLP_ECC_REG_ECC_SIGN_S_3                                                                    (32'h1000838c)
`define CLP_ECC_REG_ECC_SIGN_S_4                                                                    (32'h10008390)
`define CLP_ECC_REG_ECC_SIGN_S_5                                                                    (32'h10008394)
`define CLP_ECC_REG_ECC_SIGN_S_6                                                                    (32'h10008398)
`define CLP_ECC_REG_ECC_SIGN_S_7                                                                    (32'h1000839c)
`define CLP_ECC_REG_ECC_SIGN_S_8                                                                    (32'h100083a0)
`define CLP_ECC_REG_ECC_SIGN_S_9                                                                    (32'h100083a4)
`define CLP_ECC_REG_ECC_SIGN_S_10                                                                   (32'h100083a8)
`define CLP_ECC_REG_ECC_SIGN_S_11                                                                   (32'h100083ac)
`define CLP_ECC_REG_ECC_VERIFY_R_0                                                                  (32'h10008400)
`define CLP_ECC_REG_ECC_VERIFY_R_1                                                                  (32'h10008404)
`define CLP_ECC_REG_ECC_VERIFY_R_2                                                                  (32'h10008408)
`define CLP_ECC_REG_ECC_VERIFY_R_3                                                                  (32'h1000840c)
`define CLP_ECC_REG_ECC_VERIFY_R_4                                                                  (32'h10008410)
`define CLP_ECC_REG_ECC_VERIFY_R_5                                                                  (32'h10008414)
`define CLP_ECC_REG_ECC_VERIFY_R_6                                                                  (32'h10008418)
`define CLP_ECC_REG_ECC_VERIFY_R_7                                                                  (32'h1000841c)
`define CLP_ECC_REG_ECC_VERIFY_R_8                                                                  (32'h10008420)
`define CLP_ECC_REG_ECC_VERIFY_R_9                                                                  (32'h10008424)
`define CLP_ECC_REG_ECC_VERIFY_R_10                                                                 (32'h10008428)
`define CLP_ECC_REG_ECC_VERIFY_R_11                                                                 (32'h1000842c)
`define CLP_ECC_REG_ECC_IV_0                                                                        (32'h10008480)
`define CLP_ECC_REG_ECC_IV_1                                                                        (32'h10008484)
`define CLP_ECC_REG_ECC_IV_2                                                                        (32'h10008488)
`define CLP_ECC_REG_ECC_IV_3                                                                        (32'h1000848c)
`define CLP_ECC_REG_ECC_IV_4                                                                        (32'h10008490)
`define CLP_ECC_REG_ECC_IV_5                                                                        (32'h10008494)
`define CLP_ECC_REG_ECC_IV_6                                                                        (32'h10008498)
`define CLP_ECC_REG_ECC_IV_7                                                                        (32'h1000849c)
`define CLP_ECC_REG_ECC_IV_8                                                                        (32'h100084a0)
`define CLP_ECC_REG_ECC_IV_9                                                                        (32'h100084a4)
`define CLP_ECC_REG_ECC_IV_10                                                                       (32'h100084a8)
`define CLP_ECC_REG_ECC_IV_11                                                                       (32'h100084ac)
`define CLP_ECC_REG_ECC_NONCE_0                                                                     (32'h10008500)
`define CLP_ECC_REG_ECC_NONCE_1                                                                     (32'h10008504)
`define CLP_ECC_REG_ECC_NONCE_2                                                                     (32'h10008508)
`define CLP_ECC_REG_ECC_NONCE_3                                                                     (32'h1000850c)
`define CLP_ECC_REG_ECC_NONCE_4                                                                     (32'h10008510)
`define CLP_ECC_REG_ECC_NONCE_5                                                                     (32'h10008514)
`define CLP_ECC_REG_ECC_NONCE_6                                                                     (32'h10008518)
`define CLP_ECC_REG_ECC_NONCE_7                                                                     (32'h1000851c)
`define CLP_ECC_REG_ECC_NONCE_8                                                                     (32'h10008520)
`define CLP_ECC_REG_ECC_NONCE_9                                                                     (32'h10008524)
`define CLP_ECC_REG_ECC_NONCE_10                                                                    (32'h10008528)
`define CLP_ECC_REG_ECC_NONCE_11                                                                    (32'h1000852c)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_0                                                                (32'h10008580)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_1                                                                (32'h10008584)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_2                                                                (32'h10008588)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_3                                                                (32'h1000858c)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_4                                                                (32'h10008590)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_5                                                                (32'h10008594)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_6                                                                (32'h10008598)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_7                                                                (32'h1000859c)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_8                                                                (32'h100085a0)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_9                                                                (32'h100085a4)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_10                                                               (32'h100085a8)
`define CLP_ECC_REG_ECC_PRIVKEY_IN_11                                                               (32'h100085ac)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_0                                                             (32'h100085c0)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_1                                                             (32'h100085c4)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_2                                                             (32'h100085c8)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_3                                                             (32'h100085cc)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_4                                                             (32'h100085d0)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_5                                                             (32'h100085d4)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_6                                                             (32'h100085d8)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_7                                                             (32'h100085dc)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_8                                                             (32'h100085e0)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_9                                                             (32'h100085e4)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_10                                                            (32'h100085e8)
`define CLP_ECC_REG_ECC_DH_SHARED_KEY_11                                                            (32'h100085ec)
`define CLP_ECC_REG_ECC_KV_RD_PKEY_CTRL                                                             (32'h10008600)
`define CLP_ECC_REG_ECC_KV_RD_PKEY_STATUS                                                           (32'h10008604)
`define CLP_ECC_REG_ECC_KV_RD_SEED_CTRL                                                             (32'h10008608)
`define CLP_ECC_REG_ECC_KV_RD_SEED_STATUS                                                           (32'h1000860c)
`define CLP_ECC_REG_ECC_KV_WR_PKEY_CTRL                                                             (32'h10008610)
`define CLP_ECC_REG_ECC_KV_WR_PKEY_STATUS                                                           (32'h10008614)
`define CLP_ECC_REG_INTR_BLOCK_RF_START                                                             (32'h10008800)
`define CLP_ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10008800)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10008804)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10008808)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1000880c)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10008810)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10008814)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10008818)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1000881c)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10008820)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h10008900)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10008980)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'h10008a00)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10008a04)
`define CLP_HMAC_REG_BASE_ADDR                                                                      (32'h10010000)
`define CLP_HMAC_REG_HMAC512_NAME_0                                                                 (32'h10010000)
`define CLP_HMAC_REG_HMAC512_NAME_1                                                                 (32'h10010004)
`define CLP_HMAC_REG_HMAC512_VERSION_0                                                              (32'h10010008)
`define CLP_HMAC_REG_HMAC512_VERSION_1                                                              (32'h1001000c)
`define CLP_HMAC_REG_HMAC512_CTRL                                                                   (32'h10010010)
`define CLP_HMAC_REG_HMAC512_STATUS                                                                 (32'h10010018)
`define CLP_HMAC_REG_HMAC512_KEY_0                                                                  (32'h10010040)
`define CLP_HMAC_REG_HMAC512_KEY_1                                                                  (32'h10010044)
`define CLP_HMAC_REG_HMAC512_KEY_2                                                                  (32'h10010048)
`define CLP_HMAC_REG_HMAC512_KEY_3                                                                  (32'h1001004c)
`define CLP_HMAC_REG_HMAC512_KEY_4                                                                  (32'h10010050)
`define CLP_HMAC_REG_HMAC512_KEY_5                                                                  (32'h10010054)
`define CLP_HMAC_REG_HMAC512_KEY_6                                                                  (32'h10010058)
`define CLP_HMAC_REG_HMAC512_KEY_7                                                                  (32'h1001005c)
`define CLP_HMAC_REG_HMAC512_KEY_8                                                                  (32'h10010060)
`define CLP_HMAC_REG_HMAC512_KEY_9                                                                  (32'h10010064)
`define CLP_HMAC_REG_HMAC512_KEY_10                                                                 (32'h10010068)
`define CLP_HMAC_REG_HMAC512_KEY_11                                                                 (32'h1001006c)
`define CLP_HMAC_REG_HMAC512_KEY_12                                                                 (32'h10010070)
`define CLP_HMAC_REG_HMAC512_KEY_13                                                                 (32'h10010074)
`define CLP_HMAC_REG_HMAC512_KEY_14                                                                 (32'h10010078)
`define CLP_HMAC_REG_HMAC512_KEY_15                                                                 (32'h1001007c)
`define CLP_HMAC_REG_HMAC512_BLOCK_0                                                                (32'h10010080)
`define CLP_HMAC_REG_HMAC512_BLOCK_1                                                                (32'h10010084)
`define CLP_HMAC_REG_HMAC512_BLOCK_2                                                                (32'h10010088)
`define CLP_HMAC_REG_HMAC512_BLOCK_3                                                                (32'h1001008c)
`define CLP_HMAC_REG_HMAC512_BLOCK_4                                                                (32'h10010090)
`define CLP_HMAC_REG_HMAC512_BLOCK_5                                                                (32'h10010094)
`define CLP_HMAC_REG_HMAC512_BLOCK_6                                                                (32'h10010098)
`define CLP_HMAC_REG_HMAC512_BLOCK_7                                                                (32'h1001009c)
`define CLP_HMAC_REG_HMAC512_BLOCK_8                                                                (32'h100100a0)
`define CLP_HMAC_REG_HMAC512_BLOCK_9                                                                (32'h100100a4)
`define CLP_HMAC_REG_HMAC512_BLOCK_10                                                               (32'h100100a8)
`define CLP_HMAC_REG_HMAC512_BLOCK_11                                                               (32'h100100ac)
`define CLP_HMAC_REG_HMAC512_BLOCK_12                                                               (32'h100100b0)
`define CLP_HMAC_REG_HMAC512_BLOCK_13                                                               (32'h100100b4)
`define CLP_HMAC_REG_HMAC512_BLOCK_14                                                               (32'h100100b8)
`define CLP_HMAC_REG_HMAC512_BLOCK_15                                                               (32'h100100bc)
`define CLP_HMAC_REG_HMAC512_BLOCK_16                                                               (32'h100100c0)
`define CLP_HMAC_REG_HMAC512_BLOCK_17                                                               (32'h100100c4)
`define CLP_HMAC_REG_HMAC512_BLOCK_18                                                               (32'h100100c8)
`define CLP_HMAC_REG_HMAC512_BLOCK_19                                                               (32'h100100cc)
`define CLP_HMAC_REG_HMAC512_BLOCK_20                                                               (32'h100100d0)
`define CLP_HMAC_REG_HMAC512_BLOCK_21                                                               (32'h100100d4)
`define CLP_HMAC_REG_HMAC512_BLOCK_22                                                               (32'h100100d8)
`define CLP_HMAC_REG_HMAC512_BLOCK_23                                                               (32'h100100dc)
`define CLP_HMAC_REG_HMAC512_BLOCK_24                                                               (32'h100100e0)
`define CLP_HMAC_REG_HMAC512_BLOCK_25                                                               (32'h100100e4)
`define CLP_HMAC_REG_HMAC512_BLOCK_26                                                               (32'h100100e8)
`define CLP_HMAC_REG_HMAC512_BLOCK_27                                                               (32'h100100ec)
`define CLP_HMAC_REG_HMAC512_BLOCK_28                                                               (32'h100100f0)
`define CLP_HMAC_REG_HMAC512_BLOCK_29                                                               (32'h100100f4)
`define CLP_HMAC_REG_HMAC512_BLOCK_30                                                               (32'h100100f8)
`define CLP_HMAC_REG_HMAC512_BLOCK_31                                                               (32'h100100fc)
`define CLP_HMAC_REG_HMAC512_TAG_0                                                                  (32'h10010100)
`define CLP_HMAC_REG_HMAC512_TAG_1                                                                  (32'h10010104)
`define CLP_HMAC_REG_HMAC512_TAG_2                                                                  (32'h10010108)
`define CLP_HMAC_REG_HMAC512_TAG_3                                                                  (32'h1001010c)
`define CLP_HMAC_REG_HMAC512_TAG_4                                                                  (32'h10010110)
`define CLP_HMAC_REG_HMAC512_TAG_5                                                                  (32'h10010114)
`define CLP_HMAC_REG_HMAC512_TAG_6                                                                  (32'h10010118)
`define CLP_HMAC_REG_HMAC512_TAG_7                                                                  (32'h1001011c)
`define CLP_HMAC_REG_HMAC512_TAG_8                                                                  (32'h10010120)
`define CLP_HMAC_REG_HMAC512_TAG_9                                                                  (32'h10010124)
`define CLP_HMAC_REG_HMAC512_TAG_10                                                                 (32'h10010128)
`define CLP_HMAC_REG_HMAC512_TAG_11                                                                 (32'h1001012c)
`define CLP_HMAC_REG_HMAC512_TAG_12                                                                 (32'h10010130)
`define CLP_HMAC_REG_HMAC512_TAG_13                                                                 (32'h10010134)
`define CLP_HMAC_REG_HMAC512_TAG_14                                                                 (32'h10010138)
`define CLP_HMAC_REG_HMAC512_TAG_15                                                                 (32'h1001013c)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_0                                                            (32'h10010140)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_1                                                            (32'h10010144)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_2                                                            (32'h10010148)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_3                                                            (32'h1001014c)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_4                                                            (32'h10010150)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_5                                                            (32'h10010154)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_6                                                            (32'h10010158)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_7                                                            (32'h1001015c)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_8                                                            (32'h10010160)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_9                                                            (32'h10010164)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_10                                                           (32'h10010168)
`define CLP_HMAC_REG_HMAC512_LFSR_SEED_11                                                           (32'h1001016c)
`define CLP_HMAC_REG_HMAC512_KV_RD_KEY_CTRL                                                         (32'h10010600)
`define CLP_HMAC_REG_HMAC512_KV_RD_KEY_STATUS                                                       (32'h10010604)
`define CLP_HMAC_REG_HMAC512_KV_RD_BLOCK_CTRL                                                       (32'h10010608)
`define CLP_HMAC_REG_HMAC512_KV_RD_BLOCK_STATUS                                                     (32'h1001060c)
`define CLP_HMAC_REG_HMAC512_KV_WR_CTRL                                                             (32'h10010610)
`define CLP_HMAC_REG_HMAC512_KV_WR_STATUS                                                           (32'h10010614)
`define CLP_HMAC_REG_INTR_BLOCK_RF_START                                                            (32'h10010800)
`define CLP_HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                 (32'h10010800)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                  (32'h10010804)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                  (32'h10010808)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                              (32'h1001080c)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                              (32'h10010810)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                            (32'h10010814)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                            (32'h10010818)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                (32'h1001081c)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                (32'h10010820)
`define CLP_HMAC_REG_INTR_BLOCK_RF_KEY_MODE_ERROR_INTR_COUNT_R                                      (32'h10010900)
`define CLP_HMAC_REG_INTR_BLOCK_RF_KEY_ZERO_ERROR_INTR_COUNT_R                                      (32'h10010904)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                              (32'h10010908)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                              (32'h1001090c)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                      (32'h10010980)
`define CLP_HMAC_REG_INTR_BLOCK_RF_KEY_MODE_ERROR_INTR_COUNT_INCR_R                                 (32'h10010a00)
`define CLP_HMAC_REG_INTR_BLOCK_RF_KEY_ZERO_ERROR_INTR_COUNT_INCR_R                                 (32'h10010a04)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                         (32'h10010a08)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                         (32'h10010a0c)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                 (32'h10010a10)
`define CLP_AES_REG_BASE_ADDR                                                                       (32'h10011000)
`define CLP_AES_REG_KEY_SHARE0_0                                                                    (32'h10011004)
`define CLP_AES_REG_KEY_SHARE0_1                                                                    (32'h10011008)
`define CLP_AES_REG_KEY_SHARE0_2                                                                    (32'h1001100c)
`define CLP_AES_REG_KEY_SHARE0_3                                                                    (32'h10011010)
`define CLP_AES_REG_KEY_SHARE0_4                                                                    (32'h10011014)
`define CLP_AES_REG_KEY_SHARE0_5                                                                    (32'h10011018)
`define CLP_AES_REG_KEY_SHARE0_6                                                                    (32'h1001101c)
`define CLP_AES_REG_KEY_SHARE0_7                                                                    (32'h10011020)
`define CLP_AES_REG_KEY_SHARE1_0                                                                    (32'h10011024)
`define CLP_AES_REG_KEY_SHARE1_1                                                                    (32'h10011028)
`define CLP_AES_REG_KEY_SHARE1_2                                                                    (32'h1001102c)
`define CLP_AES_REG_KEY_SHARE1_3                                                                    (32'h10011030)
`define CLP_AES_REG_KEY_SHARE1_4                                                                    (32'h10011034)
`define CLP_AES_REG_KEY_SHARE1_5                                                                    (32'h10011038)
`define CLP_AES_REG_KEY_SHARE1_6                                                                    (32'h1001103c)
`define CLP_AES_REG_KEY_SHARE1_7                                                                    (32'h10011040)
`define CLP_AES_REG_IV_0                                                                            (32'h10011044)
`define CLP_AES_REG_IV_1                                                                            (32'h10011048)
`define CLP_AES_REG_IV_2                                                                            (32'h1001104c)
`define CLP_AES_REG_IV_3                                                                            (32'h10011050)
`define CLP_AES_REG_DATA_IN_0                                                                       (32'h10011054)
`define CLP_AES_REG_DATA_IN_1                                                                       (32'h10011058)
`define CLP_AES_REG_DATA_IN_2                                                                       (32'h1001105c)
`define CLP_AES_REG_DATA_IN_3                                                                       (32'h10011060)
`define CLP_AES_REG_DATA_OUT_0                                                                      (32'h10011064)
`define CLP_AES_REG_DATA_OUT_1                                                                      (32'h10011068)
`define CLP_AES_REG_DATA_OUT_2                                                                      (32'h1001106c)
`define CLP_AES_REG_DATA_OUT_3                                                                      (32'h10011070)
`define CLP_AES_REG_CTRL_SHADOWED                                                                   (32'h10011074)
`define CLP_AES_REG_CTRL_AUX_SHADOWED                                                               (32'h10011078)
`define CLP_AES_REG_CTRL_AUX_REGWEN                                                                 (32'h1001107c)
`define CLP_AES_REG_TRIGGER                                                                         (32'h10011080)
`define CLP_AES_REG_STATUS                                                                          (32'h10011084)
`define CLP_AES_REG_CTRL_GCM_SHADOWED                                                               (32'h10011088)
`define CLP_AES_CLP_REG_BASE_ADDR                                                                   (32'h10011800)
`define CLP_AES_CLP_REG_AES_NAME_0                                                                  (32'h10011800)
`define CLP_AES_CLP_REG_AES_NAME_1                                                                  (32'h10011804)
`define CLP_AES_CLP_REG_AES_VERSION_0                                                               (32'h10011808)
`define CLP_AES_CLP_REG_AES_VERSION_1                                                               (32'h1001180c)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_0                                                           (32'h10011910)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_1                                                           (32'h10011914)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_2                                                           (32'h10011918)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_3                                                           (32'h1001191c)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_4                                                           (32'h10011920)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_5                                                           (32'h10011924)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_6                                                           (32'h10011928)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_7                                                           (32'h1001192c)
`define CLP_AES_CLP_REG_ENTROPY_IF_SEED_8                                                           (32'h10011930)
`define CLP_AES_CLP_REG_CTRL0                                                                       (32'h10011934)
`define CLP_AES_CLP_REG_AES_KV_RD_KEY_CTRL                                                          (32'h10011a00)
`define CLP_AES_CLP_REG_AES_KV_RD_KEY_STATUS                                                        (32'h10011a04)
`define CLP_AES_CLP_REG_AES_KV_WR_CTRL                                                              (32'h10011a08)
`define CLP_AES_CLP_REG_AES_KV_WR_STATUS                                                            (32'h10011a0c)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_START                                                         (32'h10011c00)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                              (32'h10011c00)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                               (32'h10011c04)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                               (32'h10011c08)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                           (32'h10011c0c)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                           (32'h10011c10)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                         (32'h10011c14)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                         (32'h10011c18)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                             (32'h10011c1c)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                             (32'h10011c20)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                           (32'h10011d00)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                           (32'h10011d04)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                           (32'h10011d08)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                           (32'h10011d0c)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                   (32'h10011d80)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                      (32'h10011e00)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                      (32'h10011e04)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                      (32'h10011e08)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                      (32'h10011e0c)
`define CLP_AES_CLP_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                              (32'h10011e10)
`define CLP_KV_REG_BASE_ADDR                                                                        (32'h10018000)
`define CLP_KV_REG_KEY_CTRL_0                                                                       (32'h10018000)
`define CLP_KV_REG_KEY_CTRL_1                                                                       (32'h10018004)
`define CLP_KV_REG_KEY_CTRL_2                                                                       (32'h10018008)
`define CLP_KV_REG_KEY_CTRL_3                                                                       (32'h1001800c)
`define CLP_KV_REG_KEY_CTRL_4                                                                       (32'h10018010)
`define CLP_KV_REG_KEY_CTRL_5                                                                       (32'h10018014)
`define CLP_KV_REG_KEY_CTRL_6                                                                       (32'h10018018)
`define CLP_KV_REG_KEY_CTRL_7                                                                       (32'h1001801c)
`define CLP_KV_REG_KEY_CTRL_8                                                                       (32'h10018020)
`define CLP_KV_REG_KEY_CTRL_9                                                                       (32'h10018024)
`define CLP_KV_REG_KEY_CTRL_10                                                                      (32'h10018028)
`define CLP_KV_REG_KEY_CTRL_11                                                                      (32'h1001802c)
`define CLP_KV_REG_KEY_CTRL_12                                                                      (32'h10018030)
`define CLP_KV_REG_KEY_CTRL_13                                                                      (32'h10018034)
`define CLP_KV_REG_KEY_CTRL_14                                                                      (32'h10018038)
`define CLP_KV_REG_KEY_CTRL_15                                                                      (32'h1001803c)
`define CLP_KV_REG_KEY_CTRL_16                                                                      (32'h10018040)
`define CLP_KV_REG_KEY_CTRL_17                                                                      (32'h10018044)
`define CLP_KV_REG_KEY_CTRL_18                                                                      (32'h10018048)
`define CLP_KV_REG_KEY_CTRL_19                                                                      (32'h1001804c)
`define CLP_KV_REG_KEY_CTRL_20                                                                      (32'h10018050)
`define CLP_KV_REG_KEY_CTRL_21                                                                      (32'h10018054)
`define CLP_KV_REG_KEY_CTRL_22                                                                      (32'h10018058)
`define CLP_KV_REG_KEY_CTRL_23                                                                      (32'h1001805c)
`define CLP_KV_REG_KEY_ENTRY_0_0                                                                    (32'h10018600)
`define CLP_KV_REG_KEY_ENTRY_0_1                                                                    (32'h10018604)
`define CLP_KV_REG_KEY_ENTRY_0_2                                                                    (32'h10018608)
`define CLP_KV_REG_KEY_ENTRY_0_3                                                                    (32'h1001860c)
`define CLP_KV_REG_KEY_ENTRY_0_4                                                                    (32'h10018610)
`define CLP_KV_REG_KEY_ENTRY_0_5                                                                    (32'h10018614)
`define CLP_KV_REG_KEY_ENTRY_0_6                                                                    (32'h10018618)
`define CLP_KV_REG_KEY_ENTRY_0_7                                                                    (32'h1001861c)
`define CLP_KV_REG_KEY_ENTRY_0_8                                                                    (32'h10018620)
`define CLP_KV_REG_KEY_ENTRY_0_9                                                                    (32'h10018624)
`define CLP_KV_REG_KEY_ENTRY_0_10                                                                   (32'h10018628)
`define CLP_KV_REG_KEY_ENTRY_0_11                                                                   (32'h1001862c)
`define CLP_KV_REG_KEY_ENTRY_0_12                                                                   (32'h10018630)
`define CLP_KV_REG_KEY_ENTRY_0_13                                                                   (32'h10018634)
`define CLP_KV_REG_KEY_ENTRY_0_14                                                                   (32'h10018638)
`define CLP_KV_REG_KEY_ENTRY_0_15                                                                   (32'h1001863c)
`define CLP_KV_REG_KEY_ENTRY_1_0                                                                    (32'h10018640)
`define CLP_KV_REG_KEY_ENTRY_1_1                                                                    (32'h10018644)
`define CLP_KV_REG_KEY_ENTRY_1_2                                                                    (32'h10018648)
`define CLP_KV_REG_KEY_ENTRY_1_3                                                                    (32'h1001864c)
`define CLP_KV_REG_KEY_ENTRY_1_4                                                                    (32'h10018650)
`define CLP_KV_REG_KEY_ENTRY_1_5                                                                    (32'h10018654)
`define CLP_KV_REG_KEY_ENTRY_1_6                                                                    (32'h10018658)
`define CLP_KV_REG_KEY_ENTRY_1_7                                                                    (32'h1001865c)
`define CLP_KV_REG_KEY_ENTRY_1_8                                                                    (32'h10018660)
`define CLP_KV_REG_KEY_ENTRY_1_9                                                                    (32'h10018664)
`define CLP_KV_REG_KEY_ENTRY_1_10                                                                   (32'h10018668)
`define CLP_KV_REG_KEY_ENTRY_1_11                                                                   (32'h1001866c)
`define CLP_KV_REG_KEY_ENTRY_1_12                                                                   (32'h10018670)
`define CLP_KV_REG_KEY_ENTRY_1_13                                                                   (32'h10018674)
`define CLP_KV_REG_KEY_ENTRY_1_14                                                                   (32'h10018678)
`define CLP_KV_REG_KEY_ENTRY_1_15                                                                   (32'h1001867c)
`define CLP_KV_REG_KEY_ENTRY_2_0                                                                    (32'h10018680)
`define CLP_KV_REG_KEY_ENTRY_2_1                                                                    (32'h10018684)
`define CLP_KV_REG_KEY_ENTRY_2_2                                                                    (32'h10018688)
`define CLP_KV_REG_KEY_ENTRY_2_3                                                                    (32'h1001868c)
`define CLP_KV_REG_KEY_ENTRY_2_4                                                                    (32'h10018690)
`define CLP_KV_REG_KEY_ENTRY_2_5                                                                    (32'h10018694)
`define CLP_KV_REG_KEY_ENTRY_2_6                                                                    (32'h10018698)
`define CLP_KV_REG_KEY_ENTRY_2_7                                                                    (32'h1001869c)
`define CLP_KV_REG_KEY_ENTRY_2_8                                                                    (32'h100186a0)
`define CLP_KV_REG_KEY_ENTRY_2_9                                                                    (32'h100186a4)
`define CLP_KV_REG_KEY_ENTRY_2_10                                                                   (32'h100186a8)
`define CLP_KV_REG_KEY_ENTRY_2_11                                                                   (32'h100186ac)
`define CLP_KV_REG_KEY_ENTRY_2_12                                                                   (32'h100186b0)
`define CLP_KV_REG_KEY_ENTRY_2_13                                                                   (32'h100186b4)
`define CLP_KV_REG_KEY_ENTRY_2_14                                                                   (32'h100186b8)
`define CLP_KV_REG_KEY_ENTRY_2_15                                                                   (32'h100186bc)
`define CLP_KV_REG_KEY_ENTRY_3_0                                                                    (32'h100186c0)
`define CLP_KV_REG_KEY_ENTRY_3_1                                                                    (32'h100186c4)
`define CLP_KV_REG_KEY_ENTRY_3_2                                                                    (32'h100186c8)
`define CLP_KV_REG_KEY_ENTRY_3_3                                                                    (32'h100186cc)
`define CLP_KV_REG_KEY_ENTRY_3_4                                                                    (32'h100186d0)
`define CLP_KV_REG_KEY_ENTRY_3_5                                                                    (32'h100186d4)
`define CLP_KV_REG_KEY_ENTRY_3_6                                                                    (32'h100186d8)
`define CLP_KV_REG_KEY_ENTRY_3_7                                                                    (32'h100186dc)
`define CLP_KV_REG_KEY_ENTRY_3_8                                                                    (32'h100186e0)
`define CLP_KV_REG_KEY_ENTRY_3_9                                                                    (32'h100186e4)
`define CLP_KV_REG_KEY_ENTRY_3_10                                                                   (32'h100186e8)
`define CLP_KV_REG_KEY_ENTRY_3_11                                                                   (32'h100186ec)
`define CLP_KV_REG_KEY_ENTRY_3_12                                                                   (32'h100186f0)
`define CLP_KV_REG_KEY_ENTRY_3_13                                                                   (32'h100186f4)
`define CLP_KV_REG_KEY_ENTRY_3_14                                                                   (32'h100186f8)
`define CLP_KV_REG_KEY_ENTRY_3_15                                                                   (32'h100186fc)
`define CLP_KV_REG_KEY_ENTRY_4_0                                                                    (32'h10018700)
`define CLP_KV_REG_KEY_ENTRY_4_1                                                                    (32'h10018704)
`define CLP_KV_REG_KEY_ENTRY_4_2                                                                    (32'h10018708)
`define CLP_KV_REG_KEY_ENTRY_4_3                                                                    (32'h1001870c)
`define CLP_KV_REG_KEY_ENTRY_4_4                                                                    (32'h10018710)
`define CLP_KV_REG_KEY_ENTRY_4_5                                                                    (32'h10018714)
`define CLP_KV_REG_KEY_ENTRY_4_6                                                                    (32'h10018718)
`define CLP_KV_REG_KEY_ENTRY_4_7                                                                    (32'h1001871c)
`define CLP_KV_REG_KEY_ENTRY_4_8                                                                    (32'h10018720)
`define CLP_KV_REG_KEY_ENTRY_4_9                                                                    (32'h10018724)
`define CLP_KV_REG_KEY_ENTRY_4_10                                                                   (32'h10018728)
`define CLP_KV_REG_KEY_ENTRY_4_11                                                                   (32'h1001872c)
`define CLP_KV_REG_KEY_ENTRY_4_12                                                                   (32'h10018730)
`define CLP_KV_REG_KEY_ENTRY_4_13                                                                   (32'h10018734)
`define CLP_KV_REG_KEY_ENTRY_4_14                                                                   (32'h10018738)
`define CLP_KV_REG_KEY_ENTRY_4_15                                                                   (32'h1001873c)
`define CLP_KV_REG_KEY_ENTRY_5_0                                                                    (32'h10018740)
`define CLP_KV_REG_KEY_ENTRY_5_1                                                                    (32'h10018744)
`define CLP_KV_REG_KEY_ENTRY_5_2                                                                    (32'h10018748)
`define CLP_KV_REG_KEY_ENTRY_5_3                                                                    (32'h1001874c)
`define CLP_KV_REG_KEY_ENTRY_5_4                                                                    (32'h10018750)
`define CLP_KV_REG_KEY_ENTRY_5_5                                                                    (32'h10018754)
`define CLP_KV_REG_KEY_ENTRY_5_6                                                                    (32'h10018758)
`define CLP_KV_REG_KEY_ENTRY_5_7                                                                    (32'h1001875c)
`define CLP_KV_REG_KEY_ENTRY_5_8                                                                    (32'h10018760)
`define CLP_KV_REG_KEY_ENTRY_5_9                                                                    (32'h10018764)
`define CLP_KV_REG_KEY_ENTRY_5_10                                                                   (32'h10018768)
`define CLP_KV_REG_KEY_ENTRY_5_11                                                                   (32'h1001876c)
`define CLP_KV_REG_KEY_ENTRY_5_12                                                                   (32'h10018770)
`define CLP_KV_REG_KEY_ENTRY_5_13                                                                   (32'h10018774)
`define CLP_KV_REG_KEY_ENTRY_5_14                                                                   (32'h10018778)
`define CLP_KV_REG_KEY_ENTRY_5_15                                                                   (32'h1001877c)
`define CLP_KV_REG_KEY_ENTRY_6_0                                                                    (32'h10018780)
`define CLP_KV_REG_KEY_ENTRY_6_1                                                                    (32'h10018784)
`define CLP_KV_REG_KEY_ENTRY_6_2                                                                    (32'h10018788)
`define CLP_KV_REG_KEY_ENTRY_6_3                                                                    (32'h1001878c)
`define CLP_KV_REG_KEY_ENTRY_6_4                                                                    (32'h10018790)
`define CLP_KV_REG_KEY_ENTRY_6_5                                                                    (32'h10018794)
`define CLP_KV_REG_KEY_ENTRY_6_6                                                                    (32'h10018798)
`define CLP_KV_REG_KEY_ENTRY_6_7                                                                    (32'h1001879c)
`define CLP_KV_REG_KEY_ENTRY_6_8                                                                    (32'h100187a0)
`define CLP_KV_REG_KEY_ENTRY_6_9                                                                    (32'h100187a4)
`define CLP_KV_REG_KEY_ENTRY_6_10                                                                   (32'h100187a8)
`define CLP_KV_REG_KEY_ENTRY_6_11                                                                   (32'h100187ac)
`define CLP_KV_REG_KEY_ENTRY_6_12                                                                   (32'h100187b0)
`define CLP_KV_REG_KEY_ENTRY_6_13                                                                   (32'h100187b4)
`define CLP_KV_REG_KEY_ENTRY_6_14                                                                   (32'h100187b8)
`define CLP_KV_REG_KEY_ENTRY_6_15                                                                   (32'h100187bc)
`define CLP_KV_REG_KEY_ENTRY_7_0                                                                    (32'h100187c0)
`define CLP_KV_REG_KEY_ENTRY_7_1                                                                    (32'h100187c4)
`define CLP_KV_REG_KEY_ENTRY_7_2                                                                    (32'h100187c8)
`define CLP_KV_REG_KEY_ENTRY_7_3                                                                    (32'h100187cc)
`define CLP_KV_REG_KEY_ENTRY_7_4                                                                    (32'h100187d0)
`define CLP_KV_REG_KEY_ENTRY_7_5                                                                    (32'h100187d4)
`define CLP_KV_REG_KEY_ENTRY_7_6                                                                    (32'h100187d8)
`define CLP_KV_REG_KEY_ENTRY_7_7                                                                    (32'h100187dc)
`define CLP_KV_REG_KEY_ENTRY_7_8                                                                    (32'h100187e0)
`define CLP_KV_REG_KEY_ENTRY_7_9                                                                    (32'h100187e4)
`define CLP_KV_REG_KEY_ENTRY_7_10                                                                   (32'h100187e8)
`define CLP_KV_REG_KEY_ENTRY_7_11                                                                   (32'h100187ec)
`define CLP_KV_REG_KEY_ENTRY_7_12                                                                   (32'h100187f0)
`define CLP_KV_REG_KEY_ENTRY_7_13                                                                   (32'h100187f4)
`define CLP_KV_REG_KEY_ENTRY_7_14                                                                   (32'h100187f8)
`define CLP_KV_REG_KEY_ENTRY_7_15                                                                   (32'h100187fc)
`define CLP_KV_REG_KEY_ENTRY_8_0                                                                    (32'h10018800)
`define CLP_KV_REG_KEY_ENTRY_8_1                                                                    (32'h10018804)
`define CLP_KV_REG_KEY_ENTRY_8_2                                                                    (32'h10018808)
`define CLP_KV_REG_KEY_ENTRY_8_3                                                                    (32'h1001880c)
`define CLP_KV_REG_KEY_ENTRY_8_4                                                                    (32'h10018810)
`define CLP_KV_REG_KEY_ENTRY_8_5                                                                    (32'h10018814)
`define CLP_KV_REG_KEY_ENTRY_8_6                                                                    (32'h10018818)
`define CLP_KV_REG_KEY_ENTRY_8_7                                                                    (32'h1001881c)
`define CLP_KV_REG_KEY_ENTRY_8_8                                                                    (32'h10018820)
`define CLP_KV_REG_KEY_ENTRY_8_9                                                                    (32'h10018824)
`define CLP_KV_REG_KEY_ENTRY_8_10                                                                   (32'h10018828)
`define CLP_KV_REG_KEY_ENTRY_8_11                                                                   (32'h1001882c)
`define CLP_KV_REG_KEY_ENTRY_8_12                                                                   (32'h10018830)
`define CLP_KV_REG_KEY_ENTRY_8_13                                                                   (32'h10018834)
`define CLP_KV_REG_KEY_ENTRY_8_14                                                                   (32'h10018838)
`define CLP_KV_REG_KEY_ENTRY_8_15                                                                   (32'h1001883c)
`define CLP_KV_REG_KEY_ENTRY_9_0                                                                    (32'h10018840)
`define CLP_KV_REG_KEY_ENTRY_9_1                                                                    (32'h10018844)
`define CLP_KV_REG_KEY_ENTRY_9_2                                                                    (32'h10018848)
`define CLP_KV_REG_KEY_ENTRY_9_3                                                                    (32'h1001884c)
`define CLP_KV_REG_KEY_ENTRY_9_4                                                                    (32'h10018850)
`define CLP_KV_REG_KEY_ENTRY_9_5                                                                    (32'h10018854)
`define CLP_KV_REG_KEY_ENTRY_9_6                                                                    (32'h10018858)
`define CLP_KV_REG_KEY_ENTRY_9_7                                                                    (32'h1001885c)
`define CLP_KV_REG_KEY_ENTRY_9_8                                                                    (32'h10018860)
`define CLP_KV_REG_KEY_ENTRY_9_9                                                                    (32'h10018864)
`define CLP_KV_REG_KEY_ENTRY_9_10                                                                   (32'h10018868)
`define CLP_KV_REG_KEY_ENTRY_9_11                                                                   (32'h1001886c)
`define CLP_KV_REG_KEY_ENTRY_9_12                                                                   (32'h10018870)
`define CLP_KV_REG_KEY_ENTRY_9_13                                                                   (32'h10018874)
`define CLP_KV_REG_KEY_ENTRY_9_14                                                                   (32'h10018878)
`define CLP_KV_REG_KEY_ENTRY_9_15                                                                   (32'h1001887c)
`define CLP_KV_REG_KEY_ENTRY_10_0                                                                   (32'h10018880)
`define CLP_KV_REG_KEY_ENTRY_10_1                                                                   (32'h10018884)
`define CLP_KV_REG_KEY_ENTRY_10_2                                                                   (32'h10018888)
`define CLP_KV_REG_KEY_ENTRY_10_3                                                                   (32'h1001888c)
`define CLP_KV_REG_KEY_ENTRY_10_4                                                                   (32'h10018890)
`define CLP_KV_REG_KEY_ENTRY_10_5                                                                   (32'h10018894)
`define CLP_KV_REG_KEY_ENTRY_10_6                                                                   (32'h10018898)
`define CLP_KV_REG_KEY_ENTRY_10_7                                                                   (32'h1001889c)
`define CLP_KV_REG_KEY_ENTRY_10_8                                                                   (32'h100188a0)
`define CLP_KV_REG_KEY_ENTRY_10_9                                                                   (32'h100188a4)
`define CLP_KV_REG_KEY_ENTRY_10_10                                                                  (32'h100188a8)
`define CLP_KV_REG_KEY_ENTRY_10_11                                                                  (32'h100188ac)
`define CLP_KV_REG_KEY_ENTRY_10_12                                                                  (32'h100188b0)
`define CLP_KV_REG_KEY_ENTRY_10_13                                                                  (32'h100188b4)
`define CLP_KV_REG_KEY_ENTRY_10_14                                                                  (32'h100188b8)
`define CLP_KV_REG_KEY_ENTRY_10_15                                                                  (32'h100188bc)
`define CLP_KV_REG_KEY_ENTRY_11_0                                                                   (32'h100188c0)
`define CLP_KV_REG_KEY_ENTRY_11_1                                                                   (32'h100188c4)
`define CLP_KV_REG_KEY_ENTRY_11_2                                                                   (32'h100188c8)
`define CLP_KV_REG_KEY_ENTRY_11_3                                                                   (32'h100188cc)
`define CLP_KV_REG_KEY_ENTRY_11_4                                                                   (32'h100188d0)
`define CLP_KV_REG_KEY_ENTRY_11_5                                                                   (32'h100188d4)
`define CLP_KV_REG_KEY_ENTRY_11_6                                                                   (32'h100188d8)
`define CLP_KV_REG_KEY_ENTRY_11_7                                                                   (32'h100188dc)
`define CLP_KV_REG_KEY_ENTRY_11_8                                                                   (32'h100188e0)
`define CLP_KV_REG_KEY_ENTRY_11_9                                                                   (32'h100188e4)
`define CLP_KV_REG_KEY_ENTRY_11_10                                                                  (32'h100188e8)
`define CLP_KV_REG_KEY_ENTRY_11_11                                                                  (32'h100188ec)
`define CLP_KV_REG_KEY_ENTRY_11_12                                                                  (32'h100188f0)
`define CLP_KV_REG_KEY_ENTRY_11_13                                                                  (32'h100188f4)
`define CLP_KV_REG_KEY_ENTRY_11_14                                                                  (32'h100188f8)
`define CLP_KV_REG_KEY_ENTRY_11_15                                                                  (32'h100188fc)
`define CLP_KV_REG_KEY_ENTRY_12_0                                                                   (32'h10018900)
`define CLP_KV_REG_KEY_ENTRY_12_1                                                                   (32'h10018904)
`define CLP_KV_REG_KEY_ENTRY_12_2                                                                   (32'h10018908)
`define CLP_KV_REG_KEY_ENTRY_12_3                                                                   (32'h1001890c)
`define CLP_KV_REG_KEY_ENTRY_12_4                                                                   (32'h10018910)
`define CLP_KV_REG_KEY_ENTRY_12_5                                                                   (32'h10018914)
`define CLP_KV_REG_KEY_ENTRY_12_6                                                                   (32'h10018918)
`define CLP_KV_REG_KEY_ENTRY_12_7                                                                   (32'h1001891c)
`define CLP_KV_REG_KEY_ENTRY_12_8                                                                   (32'h10018920)
`define CLP_KV_REG_KEY_ENTRY_12_9                                                                   (32'h10018924)
`define CLP_KV_REG_KEY_ENTRY_12_10                                                                  (32'h10018928)
`define CLP_KV_REG_KEY_ENTRY_12_11                                                                  (32'h1001892c)
`define CLP_KV_REG_KEY_ENTRY_12_12                                                                  (32'h10018930)
`define CLP_KV_REG_KEY_ENTRY_12_13                                                                  (32'h10018934)
`define CLP_KV_REG_KEY_ENTRY_12_14                                                                  (32'h10018938)
`define CLP_KV_REG_KEY_ENTRY_12_15                                                                  (32'h1001893c)
`define CLP_KV_REG_KEY_ENTRY_13_0                                                                   (32'h10018940)
`define CLP_KV_REG_KEY_ENTRY_13_1                                                                   (32'h10018944)
`define CLP_KV_REG_KEY_ENTRY_13_2                                                                   (32'h10018948)
`define CLP_KV_REG_KEY_ENTRY_13_3                                                                   (32'h1001894c)
`define CLP_KV_REG_KEY_ENTRY_13_4                                                                   (32'h10018950)
`define CLP_KV_REG_KEY_ENTRY_13_5                                                                   (32'h10018954)
`define CLP_KV_REG_KEY_ENTRY_13_6                                                                   (32'h10018958)
`define CLP_KV_REG_KEY_ENTRY_13_7                                                                   (32'h1001895c)
`define CLP_KV_REG_KEY_ENTRY_13_8                                                                   (32'h10018960)
`define CLP_KV_REG_KEY_ENTRY_13_9                                                                   (32'h10018964)
`define CLP_KV_REG_KEY_ENTRY_13_10                                                                  (32'h10018968)
`define CLP_KV_REG_KEY_ENTRY_13_11                                                                  (32'h1001896c)
`define CLP_KV_REG_KEY_ENTRY_13_12                                                                  (32'h10018970)
`define CLP_KV_REG_KEY_ENTRY_13_13                                                                  (32'h10018974)
`define CLP_KV_REG_KEY_ENTRY_13_14                                                                  (32'h10018978)
`define CLP_KV_REG_KEY_ENTRY_13_15                                                                  (32'h1001897c)
`define CLP_KV_REG_KEY_ENTRY_14_0                                                                   (32'h10018980)
`define CLP_KV_REG_KEY_ENTRY_14_1                                                                   (32'h10018984)
`define CLP_KV_REG_KEY_ENTRY_14_2                                                                   (32'h10018988)
`define CLP_KV_REG_KEY_ENTRY_14_3                                                                   (32'h1001898c)
`define CLP_KV_REG_KEY_ENTRY_14_4                                                                   (32'h10018990)
`define CLP_KV_REG_KEY_ENTRY_14_5                                                                   (32'h10018994)
`define CLP_KV_REG_KEY_ENTRY_14_6                                                                   (32'h10018998)
`define CLP_KV_REG_KEY_ENTRY_14_7                                                                   (32'h1001899c)
`define CLP_KV_REG_KEY_ENTRY_14_8                                                                   (32'h100189a0)
`define CLP_KV_REG_KEY_ENTRY_14_9                                                                   (32'h100189a4)
`define CLP_KV_REG_KEY_ENTRY_14_10                                                                  (32'h100189a8)
`define CLP_KV_REG_KEY_ENTRY_14_11                                                                  (32'h100189ac)
`define CLP_KV_REG_KEY_ENTRY_14_12                                                                  (32'h100189b0)
`define CLP_KV_REG_KEY_ENTRY_14_13                                                                  (32'h100189b4)
`define CLP_KV_REG_KEY_ENTRY_14_14                                                                  (32'h100189b8)
`define CLP_KV_REG_KEY_ENTRY_14_15                                                                  (32'h100189bc)
`define CLP_KV_REG_KEY_ENTRY_15_0                                                                   (32'h100189c0)
`define CLP_KV_REG_KEY_ENTRY_15_1                                                                   (32'h100189c4)
`define CLP_KV_REG_KEY_ENTRY_15_2                                                                   (32'h100189c8)
`define CLP_KV_REG_KEY_ENTRY_15_3                                                                   (32'h100189cc)
`define CLP_KV_REG_KEY_ENTRY_15_4                                                                   (32'h100189d0)
`define CLP_KV_REG_KEY_ENTRY_15_5                                                                   (32'h100189d4)
`define CLP_KV_REG_KEY_ENTRY_15_6                                                                   (32'h100189d8)
`define CLP_KV_REG_KEY_ENTRY_15_7                                                                   (32'h100189dc)
`define CLP_KV_REG_KEY_ENTRY_15_8                                                                   (32'h100189e0)
`define CLP_KV_REG_KEY_ENTRY_15_9                                                                   (32'h100189e4)
`define CLP_KV_REG_KEY_ENTRY_15_10                                                                  (32'h100189e8)
`define CLP_KV_REG_KEY_ENTRY_15_11                                                                  (32'h100189ec)
`define CLP_KV_REG_KEY_ENTRY_15_12                                                                  (32'h100189f0)
`define CLP_KV_REG_KEY_ENTRY_15_13                                                                  (32'h100189f4)
`define CLP_KV_REG_KEY_ENTRY_15_14                                                                  (32'h100189f8)
`define CLP_KV_REG_KEY_ENTRY_15_15                                                                  (32'h100189fc)
`define CLP_KV_REG_KEY_ENTRY_16_0                                                                   (32'h10018a00)
`define CLP_KV_REG_KEY_ENTRY_16_1                                                                   (32'h10018a04)
`define CLP_KV_REG_KEY_ENTRY_16_2                                                                   (32'h10018a08)
`define CLP_KV_REG_KEY_ENTRY_16_3                                                                   (32'h10018a0c)
`define CLP_KV_REG_KEY_ENTRY_16_4                                                                   (32'h10018a10)
`define CLP_KV_REG_KEY_ENTRY_16_5                                                                   (32'h10018a14)
`define CLP_KV_REG_KEY_ENTRY_16_6                                                                   (32'h10018a18)
`define CLP_KV_REG_KEY_ENTRY_16_7                                                                   (32'h10018a1c)
`define CLP_KV_REG_KEY_ENTRY_16_8                                                                   (32'h10018a20)
`define CLP_KV_REG_KEY_ENTRY_16_9                                                                   (32'h10018a24)
`define CLP_KV_REG_KEY_ENTRY_16_10                                                                  (32'h10018a28)
`define CLP_KV_REG_KEY_ENTRY_16_11                                                                  (32'h10018a2c)
`define CLP_KV_REG_KEY_ENTRY_16_12                                                                  (32'h10018a30)
`define CLP_KV_REG_KEY_ENTRY_16_13                                                                  (32'h10018a34)
`define CLP_KV_REG_KEY_ENTRY_16_14                                                                  (32'h10018a38)
`define CLP_KV_REG_KEY_ENTRY_16_15                                                                  (32'h10018a3c)
`define CLP_KV_REG_KEY_ENTRY_17_0                                                                   (32'h10018a40)
`define CLP_KV_REG_KEY_ENTRY_17_1                                                                   (32'h10018a44)
`define CLP_KV_REG_KEY_ENTRY_17_2                                                                   (32'h10018a48)
`define CLP_KV_REG_KEY_ENTRY_17_3                                                                   (32'h10018a4c)
`define CLP_KV_REG_KEY_ENTRY_17_4                                                                   (32'h10018a50)
`define CLP_KV_REG_KEY_ENTRY_17_5                                                                   (32'h10018a54)
`define CLP_KV_REG_KEY_ENTRY_17_6                                                                   (32'h10018a58)
`define CLP_KV_REG_KEY_ENTRY_17_7                                                                   (32'h10018a5c)
`define CLP_KV_REG_KEY_ENTRY_17_8                                                                   (32'h10018a60)
`define CLP_KV_REG_KEY_ENTRY_17_9                                                                   (32'h10018a64)
`define CLP_KV_REG_KEY_ENTRY_17_10                                                                  (32'h10018a68)
`define CLP_KV_REG_KEY_ENTRY_17_11                                                                  (32'h10018a6c)
`define CLP_KV_REG_KEY_ENTRY_17_12                                                                  (32'h10018a70)
`define CLP_KV_REG_KEY_ENTRY_17_13                                                                  (32'h10018a74)
`define CLP_KV_REG_KEY_ENTRY_17_14                                                                  (32'h10018a78)
`define CLP_KV_REG_KEY_ENTRY_17_15                                                                  (32'h10018a7c)
`define CLP_KV_REG_KEY_ENTRY_18_0                                                                   (32'h10018a80)
`define CLP_KV_REG_KEY_ENTRY_18_1                                                                   (32'h10018a84)
`define CLP_KV_REG_KEY_ENTRY_18_2                                                                   (32'h10018a88)
`define CLP_KV_REG_KEY_ENTRY_18_3                                                                   (32'h10018a8c)
`define CLP_KV_REG_KEY_ENTRY_18_4                                                                   (32'h10018a90)
`define CLP_KV_REG_KEY_ENTRY_18_5                                                                   (32'h10018a94)
`define CLP_KV_REG_KEY_ENTRY_18_6                                                                   (32'h10018a98)
`define CLP_KV_REG_KEY_ENTRY_18_7                                                                   (32'h10018a9c)
`define CLP_KV_REG_KEY_ENTRY_18_8                                                                   (32'h10018aa0)
`define CLP_KV_REG_KEY_ENTRY_18_9                                                                   (32'h10018aa4)
`define CLP_KV_REG_KEY_ENTRY_18_10                                                                  (32'h10018aa8)
`define CLP_KV_REG_KEY_ENTRY_18_11                                                                  (32'h10018aac)
`define CLP_KV_REG_KEY_ENTRY_18_12                                                                  (32'h10018ab0)
`define CLP_KV_REG_KEY_ENTRY_18_13                                                                  (32'h10018ab4)
`define CLP_KV_REG_KEY_ENTRY_18_14                                                                  (32'h10018ab8)
`define CLP_KV_REG_KEY_ENTRY_18_15                                                                  (32'h10018abc)
`define CLP_KV_REG_KEY_ENTRY_19_0                                                                   (32'h10018ac0)
`define CLP_KV_REG_KEY_ENTRY_19_1                                                                   (32'h10018ac4)
`define CLP_KV_REG_KEY_ENTRY_19_2                                                                   (32'h10018ac8)
`define CLP_KV_REG_KEY_ENTRY_19_3                                                                   (32'h10018acc)
`define CLP_KV_REG_KEY_ENTRY_19_4                                                                   (32'h10018ad0)
`define CLP_KV_REG_KEY_ENTRY_19_5                                                                   (32'h10018ad4)
`define CLP_KV_REG_KEY_ENTRY_19_6                                                                   (32'h10018ad8)
`define CLP_KV_REG_KEY_ENTRY_19_7                                                                   (32'h10018adc)
`define CLP_KV_REG_KEY_ENTRY_19_8                                                                   (32'h10018ae0)
`define CLP_KV_REG_KEY_ENTRY_19_9                                                                   (32'h10018ae4)
`define CLP_KV_REG_KEY_ENTRY_19_10                                                                  (32'h10018ae8)
`define CLP_KV_REG_KEY_ENTRY_19_11                                                                  (32'h10018aec)
`define CLP_KV_REG_KEY_ENTRY_19_12                                                                  (32'h10018af0)
`define CLP_KV_REG_KEY_ENTRY_19_13                                                                  (32'h10018af4)
`define CLP_KV_REG_KEY_ENTRY_19_14                                                                  (32'h10018af8)
`define CLP_KV_REG_KEY_ENTRY_19_15                                                                  (32'h10018afc)
`define CLP_KV_REG_KEY_ENTRY_20_0                                                                   (32'h10018b00)
`define CLP_KV_REG_KEY_ENTRY_20_1                                                                   (32'h10018b04)
`define CLP_KV_REG_KEY_ENTRY_20_2                                                                   (32'h10018b08)
`define CLP_KV_REG_KEY_ENTRY_20_3                                                                   (32'h10018b0c)
`define CLP_KV_REG_KEY_ENTRY_20_4                                                                   (32'h10018b10)
`define CLP_KV_REG_KEY_ENTRY_20_5                                                                   (32'h10018b14)
`define CLP_KV_REG_KEY_ENTRY_20_6                                                                   (32'h10018b18)
`define CLP_KV_REG_KEY_ENTRY_20_7                                                                   (32'h10018b1c)
`define CLP_KV_REG_KEY_ENTRY_20_8                                                                   (32'h10018b20)
`define CLP_KV_REG_KEY_ENTRY_20_9                                                                   (32'h10018b24)
`define CLP_KV_REG_KEY_ENTRY_20_10                                                                  (32'h10018b28)
`define CLP_KV_REG_KEY_ENTRY_20_11                                                                  (32'h10018b2c)
`define CLP_KV_REG_KEY_ENTRY_20_12                                                                  (32'h10018b30)
`define CLP_KV_REG_KEY_ENTRY_20_13                                                                  (32'h10018b34)
`define CLP_KV_REG_KEY_ENTRY_20_14                                                                  (32'h10018b38)
`define CLP_KV_REG_KEY_ENTRY_20_15                                                                  (32'h10018b3c)
`define CLP_KV_REG_KEY_ENTRY_21_0                                                                   (32'h10018b40)
`define CLP_KV_REG_KEY_ENTRY_21_1                                                                   (32'h10018b44)
`define CLP_KV_REG_KEY_ENTRY_21_2                                                                   (32'h10018b48)
`define CLP_KV_REG_KEY_ENTRY_21_3                                                                   (32'h10018b4c)
`define CLP_KV_REG_KEY_ENTRY_21_4                                                                   (32'h10018b50)
`define CLP_KV_REG_KEY_ENTRY_21_5                                                                   (32'h10018b54)
`define CLP_KV_REG_KEY_ENTRY_21_6                                                                   (32'h10018b58)
`define CLP_KV_REG_KEY_ENTRY_21_7                                                                   (32'h10018b5c)
`define CLP_KV_REG_KEY_ENTRY_21_8                                                                   (32'h10018b60)
`define CLP_KV_REG_KEY_ENTRY_21_9                                                                   (32'h10018b64)
`define CLP_KV_REG_KEY_ENTRY_21_10                                                                  (32'h10018b68)
`define CLP_KV_REG_KEY_ENTRY_21_11                                                                  (32'h10018b6c)
`define CLP_KV_REG_KEY_ENTRY_21_12                                                                  (32'h10018b70)
`define CLP_KV_REG_KEY_ENTRY_21_13                                                                  (32'h10018b74)
`define CLP_KV_REG_KEY_ENTRY_21_14                                                                  (32'h10018b78)
`define CLP_KV_REG_KEY_ENTRY_21_15                                                                  (32'h10018b7c)
`define CLP_KV_REG_KEY_ENTRY_22_0                                                                   (32'h10018b80)
`define CLP_KV_REG_KEY_ENTRY_22_1                                                                   (32'h10018b84)
`define CLP_KV_REG_KEY_ENTRY_22_2                                                                   (32'h10018b88)
`define CLP_KV_REG_KEY_ENTRY_22_3                                                                   (32'h10018b8c)
`define CLP_KV_REG_KEY_ENTRY_22_4                                                                   (32'h10018b90)
`define CLP_KV_REG_KEY_ENTRY_22_5                                                                   (32'h10018b94)
`define CLP_KV_REG_KEY_ENTRY_22_6                                                                   (32'h10018b98)
`define CLP_KV_REG_KEY_ENTRY_22_7                                                                   (32'h10018b9c)
`define CLP_KV_REG_KEY_ENTRY_22_8                                                                   (32'h10018ba0)
`define CLP_KV_REG_KEY_ENTRY_22_9                                                                   (32'h10018ba4)
`define CLP_KV_REG_KEY_ENTRY_22_10                                                                  (32'h10018ba8)
`define CLP_KV_REG_KEY_ENTRY_22_11                                                                  (32'h10018bac)
`define CLP_KV_REG_KEY_ENTRY_22_12                                                                  (32'h10018bb0)
`define CLP_KV_REG_KEY_ENTRY_22_13                                                                  (32'h10018bb4)
`define CLP_KV_REG_KEY_ENTRY_22_14                                                                  (32'h10018bb8)
`define CLP_KV_REG_KEY_ENTRY_22_15                                                                  (32'h10018bbc)
`define CLP_KV_REG_KEY_ENTRY_23_0                                                                   (32'h10018bc0)
`define CLP_KV_REG_KEY_ENTRY_23_1                                                                   (32'h10018bc4)
`define CLP_KV_REG_KEY_ENTRY_23_2                                                                   (32'h10018bc8)
`define CLP_KV_REG_KEY_ENTRY_23_3                                                                   (32'h10018bcc)
`define CLP_KV_REG_KEY_ENTRY_23_4                                                                   (32'h10018bd0)
`define CLP_KV_REG_KEY_ENTRY_23_5                                                                   (32'h10018bd4)
`define CLP_KV_REG_KEY_ENTRY_23_6                                                                   (32'h10018bd8)
`define CLP_KV_REG_KEY_ENTRY_23_7                                                                   (32'h10018bdc)
`define CLP_KV_REG_KEY_ENTRY_23_8                                                                   (32'h10018be0)
`define CLP_KV_REG_KEY_ENTRY_23_9                                                                   (32'h10018be4)
`define CLP_KV_REG_KEY_ENTRY_23_10                                                                  (32'h10018be8)
`define CLP_KV_REG_KEY_ENTRY_23_11                                                                  (32'h10018bec)
`define CLP_KV_REG_KEY_ENTRY_23_12                                                                  (32'h10018bf0)
`define CLP_KV_REG_KEY_ENTRY_23_13                                                                  (32'h10018bf4)
`define CLP_KV_REG_KEY_ENTRY_23_14                                                                  (32'h10018bf8)
`define CLP_KV_REG_KEY_ENTRY_23_15                                                                  (32'h10018bfc)
`define CLP_KV_REG_CLEAR_SECRETS                                                                    (32'h10018c00)
`define CLP_PV_REG_BASE_ADDR                                                                        (32'h1001a000)
`define CLP_PV_REG_PCR_CTRL_0                                                                       (32'h1001a000)
`define CLP_PV_REG_PCR_CTRL_1                                                                       (32'h1001a004)
`define CLP_PV_REG_PCR_CTRL_2                                                                       (32'h1001a008)
`define CLP_PV_REG_PCR_CTRL_3                                                                       (32'h1001a00c)
`define CLP_PV_REG_PCR_CTRL_4                                                                       (32'h1001a010)
`define CLP_PV_REG_PCR_CTRL_5                                                                       (32'h1001a014)
`define CLP_PV_REG_PCR_CTRL_6                                                                       (32'h1001a018)
`define CLP_PV_REG_PCR_CTRL_7                                                                       (32'h1001a01c)
`define CLP_PV_REG_PCR_CTRL_8                                                                       (32'h1001a020)
`define CLP_PV_REG_PCR_CTRL_9                                                                       (32'h1001a024)
`define CLP_PV_REG_PCR_CTRL_10                                                                      (32'h1001a028)
`define CLP_PV_REG_PCR_CTRL_11                                                                      (32'h1001a02c)
`define CLP_PV_REG_PCR_CTRL_12                                                                      (32'h1001a030)
`define CLP_PV_REG_PCR_CTRL_13                                                                      (32'h1001a034)
`define CLP_PV_REG_PCR_CTRL_14                                                                      (32'h1001a038)
`define CLP_PV_REG_PCR_CTRL_15                                                                      (32'h1001a03c)
`define CLP_PV_REG_PCR_CTRL_16                                                                      (32'h1001a040)
`define CLP_PV_REG_PCR_CTRL_17                                                                      (32'h1001a044)
`define CLP_PV_REG_PCR_CTRL_18                                                                      (32'h1001a048)
`define CLP_PV_REG_PCR_CTRL_19                                                                      (32'h1001a04c)
`define CLP_PV_REG_PCR_CTRL_20                                                                      (32'h1001a050)
`define CLP_PV_REG_PCR_CTRL_21                                                                      (32'h1001a054)
`define CLP_PV_REG_PCR_CTRL_22                                                                      (32'h1001a058)
`define CLP_PV_REG_PCR_CTRL_23                                                                      (32'h1001a05c)
`define CLP_PV_REG_PCR_CTRL_24                                                                      (32'h1001a060)
`define CLP_PV_REG_PCR_CTRL_25                                                                      (32'h1001a064)
`define CLP_PV_REG_PCR_CTRL_26                                                                      (32'h1001a068)
`define CLP_PV_REG_PCR_CTRL_27                                                                      (32'h1001a06c)
`define CLP_PV_REG_PCR_CTRL_28                                                                      (32'h1001a070)
`define CLP_PV_REG_PCR_CTRL_29                                                                      (32'h1001a074)
`define CLP_PV_REG_PCR_CTRL_30                                                                      (32'h1001a078)
`define CLP_PV_REG_PCR_CTRL_31                                                                      (32'h1001a07c)
`define CLP_PV_REG_PCR_ENTRY_0_0                                                                    (32'h1001a600)
`define CLP_PV_REG_PCR_ENTRY_0_1                                                                    (32'h1001a604)
`define CLP_PV_REG_PCR_ENTRY_0_2                                                                    (32'h1001a608)
`define CLP_PV_REG_PCR_ENTRY_0_3                                                                    (32'h1001a60c)
`define CLP_PV_REG_PCR_ENTRY_0_4                                                                    (32'h1001a610)
`define CLP_PV_REG_PCR_ENTRY_0_5                                                                    (32'h1001a614)
`define CLP_PV_REG_PCR_ENTRY_0_6                                                                    (32'h1001a618)
`define CLP_PV_REG_PCR_ENTRY_0_7                                                                    (32'h1001a61c)
`define CLP_PV_REG_PCR_ENTRY_0_8                                                                    (32'h1001a620)
`define CLP_PV_REG_PCR_ENTRY_0_9                                                                    (32'h1001a624)
`define CLP_PV_REG_PCR_ENTRY_0_10                                                                   (32'h1001a628)
`define CLP_PV_REG_PCR_ENTRY_0_11                                                                   (32'h1001a62c)
`define CLP_PV_REG_PCR_ENTRY_1_0                                                                    (32'h1001a630)
`define CLP_PV_REG_PCR_ENTRY_1_1                                                                    (32'h1001a634)
`define CLP_PV_REG_PCR_ENTRY_1_2                                                                    (32'h1001a638)
`define CLP_PV_REG_PCR_ENTRY_1_3                                                                    (32'h1001a63c)
`define CLP_PV_REG_PCR_ENTRY_1_4                                                                    (32'h1001a640)
`define CLP_PV_REG_PCR_ENTRY_1_5                                                                    (32'h1001a644)
`define CLP_PV_REG_PCR_ENTRY_1_6                                                                    (32'h1001a648)
`define CLP_PV_REG_PCR_ENTRY_1_7                                                                    (32'h1001a64c)
`define CLP_PV_REG_PCR_ENTRY_1_8                                                                    (32'h1001a650)
`define CLP_PV_REG_PCR_ENTRY_1_9                                                                    (32'h1001a654)
`define CLP_PV_REG_PCR_ENTRY_1_10                                                                   (32'h1001a658)
`define CLP_PV_REG_PCR_ENTRY_1_11                                                                   (32'h1001a65c)
`define CLP_PV_REG_PCR_ENTRY_2_0                                                                    (32'h1001a660)
`define CLP_PV_REG_PCR_ENTRY_2_1                                                                    (32'h1001a664)
`define CLP_PV_REG_PCR_ENTRY_2_2                                                                    (32'h1001a668)
`define CLP_PV_REG_PCR_ENTRY_2_3                                                                    (32'h1001a66c)
`define CLP_PV_REG_PCR_ENTRY_2_4                                                                    (32'h1001a670)
`define CLP_PV_REG_PCR_ENTRY_2_5                                                                    (32'h1001a674)
`define CLP_PV_REG_PCR_ENTRY_2_6                                                                    (32'h1001a678)
`define CLP_PV_REG_PCR_ENTRY_2_7                                                                    (32'h1001a67c)
`define CLP_PV_REG_PCR_ENTRY_2_8                                                                    (32'h1001a680)
`define CLP_PV_REG_PCR_ENTRY_2_9                                                                    (32'h1001a684)
`define CLP_PV_REG_PCR_ENTRY_2_10                                                                   (32'h1001a688)
`define CLP_PV_REG_PCR_ENTRY_2_11                                                                   (32'h1001a68c)
`define CLP_PV_REG_PCR_ENTRY_3_0                                                                    (32'h1001a690)
`define CLP_PV_REG_PCR_ENTRY_3_1                                                                    (32'h1001a694)
`define CLP_PV_REG_PCR_ENTRY_3_2                                                                    (32'h1001a698)
`define CLP_PV_REG_PCR_ENTRY_3_3                                                                    (32'h1001a69c)
`define CLP_PV_REG_PCR_ENTRY_3_4                                                                    (32'h1001a6a0)
`define CLP_PV_REG_PCR_ENTRY_3_5                                                                    (32'h1001a6a4)
`define CLP_PV_REG_PCR_ENTRY_3_6                                                                    (32'h1001a6a8)
`define CLP_PV_REG_PCR_ENTRY_3_7                                                                    (32'h1001a6ac)
`define CLP_PV_REG_PCR_ENTRY_3_8                                                                    (32'h1001a6b0)
`define CLP_PV_REG_PCR_ENTRY_3_9                                                                    (32'h1001a6b4)
`define CLP_PV_REG_PCR_ENTRY_3_10                                                                   (32'h1001a6b8)
`define CLP_PV_REG_PCR_ENTRY_3_11                                                                   (32'h1001a6bc)
`define CLP_PV_REG_PCR_ENTRY_4_0                                                                    (32'h1001a6c0)
`define CLP_PV_REG_PCR_ENTRY_4_1                                                                    (32'h1001a6c4)
`define CLP_PV_REG_PCR_ENTRY_4_2                                                                    (32'h1001a6c8)
`define CLP_PV_REG_PCR_ENTRY_4_3                                                                    (32'h1001a6cc)
`define CLP_PV_REG_PCR_ENTRY_4_4                                                                    (32'h1001a6d0)
`define CLP_PV_REG_PCR_ENTRY_4_5                                                                    (32'h1001a6d4)
`define CLP_PV_REG_PCR_ENTRY_4_6                                                                    (32'h1001a6d8)
`define CLP_PV_REG_PCR_ENTRY_4_7                                                                    (32'h1001a6dc)
`define CLP_PV_REG_PCR_ENTRY_4_8                                                                    (32'h1001a6e0)
`define CLP_PV_REG_PCR_ENTRY_4_9                                                                    (32'h1001a6e4)
`define CLP_PV_REG_PCR_ENTRY_4_10                                                                   (32'h1001a6e8)
`define CLP_PV_REG_PCR_ENTRY_4_11                                                                   (32'h1001a6ec)
`define CLP_PV_REG_PCR_ENTRY_5_0                                                                    (32'h1001a6f0)
`define CLP_PV_REG_PCR_ENTRY_5_1                                                                    (32'h1001a6f4)
`define CLP_PV_REG_PCR_ENTRY_5_2                                                                    (32'h1001a6f8)
`define CLP_PV_REG_PCR_ENTRY_5_3                                                                    (32'h1001a6fc)
`define CLP_PV_REG_PCR_ENTRY_5_4                                                                    (32'h1001a700)
`define CLP_PV_REG_PCR_ENTRY_5_5                                                                    (32'h1001a704)
`define CLP_PV_REG_PCR_ENTRY_5_6                                                                    (32'h1001a708)
`define CLP_PV_REG_PCR_ENTRY_5_7                                                                    (32'h1001a70c)
`define CLP_PV_REG_PCR_ENTRY_5_8                                                                    (32'h1001a710)
`define CLP_PV_REG_PCR_ENTRY_5_9                                                                    (32'h1001a714)
`define CLP_PV_REG_PCR_ENTRY_5_10                                                                   (32'h1001a718)
`define CLP_PV_REG_PCR_ENTRY_5_11                                                                   (32'h1001a71c)
`define CLP_PV_REG_PCR_ENTRY_6_0                                                                    (32'h1001a720)
`define CLP_PV_REG_PCR_ENTRY_6_1                                                                    (32'h1001a724)
`define CLP_PV_REG_PCR_ENTRY_6_2                                                                    (32'h1001a728)
`define CLP_PV_REG_PCR_ENTRY_6_3                                                                    (32'h1001a72c)
`define CLP_PV_REG_PCR_ENTRY_6_4                                                                    (32'h1001a730)
`define CLP_PV_REG_PCR_ENTRY_6_5                                                                    (32'h1001a734)
`define CLP_PV_REG_PCR_ENTRY_6_6                                                                    (32'h1001a738)
`define CLP_PV_REG_PCR_ENTRY_6_7                                                                    (32'h1001a73c)
`define CLP_PV_REG_PCR_ENTRY_6_8                                                                    (32'h1001a740)
`define CLP_PV_REG_PCR_ENTRY_6_9                                                                    (32'h1001a744)
`define CLP_PV_REG_PCR_ENTRY_6_10                                                                   (32'h1001a748)
`define CLP_PV_REG_PCR_ENTRY_6_11                                                                   (32'h1001a74c)
`define CLP_PV_REG_PCR_ENTRY_7_0                                                                    (32'h1001a750)
`define CLP_PV_REG_PCR_ENTRY_7_1                                                                    (32'h1001a754)
`define CLP_PV_REG_PCR_ENTRY_7_2                                                                    (32'h1001a758)
`define CLP_PV_REG_PCR_ENTRY_7_3                                                                    (32'h1001a75c)
`define CLP_PV_REG_PCR_ENTRY_7_4                                                                    (32'h1001a760)
`define CLP_PV_REG_PCR_ENTRY_7_5                                                                    (32'h1001a764)
`define CLP_PV_REG_PCR_ENTRY_7_6                                                                    (32'h1001a768)
`define CLP_PV_REG_PCR_ENTRY_7_7                                                                    (32'h1001a76c)
`define CLP_PV_REG_PCR_ENTRY_7_8                                                                    (32'h1001a770)
`define CLP_PV_REG_PCR_ENTRY_7_9                                                                    (32'h1001a774)
`define CLP_PV_REG_PCR_ENTRY_7_10                                                                   (32'h1001a778)
`define CLP_PV_REG_PCR_ENTRY_7_11                                                                   (32'h1001a77c)
`define CLP_PV_REG_PCR_ENTRY_8_0                                                                    (32'h1001a780)
`define CLP_PV_REG_PCR_ENTRY_8_1                                                                    (32'h1001a784)
`define CLP_PV_REG_PCR_ENTRY_8_2                                                                    (32'h1001a788)
`define CLP_PV_REG_PCR_ENTRY_8_3                                                                    (32'h1001a78c)
`define CLP_PV_REG_PCR_ENTRY_8_4                                                                    (32'h1001a790)
`define CLP_PV_REG_PCR_ENTRY_8_5                                                                    (32'h1001a794)
`define CLP_PV_REG_PCR_ENTRY_8_6                                                                    (32'h1001a798)
`define CLP_PV_REG_PCR_ENTRY_8_7                                                                    (32'h1001a79c)
`define CLP_PV_REG_PCR_ENTRY_8_8                                                                    (32'h1001a7a0)
`define CLP_PV_REG_PCR_ENTRY_8_9                                                                    (32'h1001a7a4)
`define CLP_PV_REG_PCR_ENTRY_8_10                                                                   (32'h1001a7a8)
`define CLP_PV_REG_PCR_ENTRY_8_11                                                                   (32'h1001a7ac)
`define CLP_PV_REG_PCR_ENTRY_9_0                                                                    (32'h1001a7b0)
`define CLP_PV_REG_PCR_ENTRY_9_1                                                                    (32'h1001a7b4)
`define CLP_PV_REG_PCR_ENTRY_9_2                                                                    (32'h1001a7b8)
`define CLP_PV_REG_PCR_ENTRY_9_3                                                                    (32'h1001a7bc)
`define CLP_PV_REG_PCR_ENTRY_9_4                                                                    (32'h1001a7c0)
`define CLP_PV_REG_PCR_ENTRY_9_5                                                                    (32'h1001a7c4)
`define CLP_PV_REG_PCR_ENTRY_9_6                                                                    (32'h1001a7c8)
`define CLP_PV_REG_PCR_ENTRY_9_7                                                                    (32'h1001a7cc)
`define CLP_PV_REG_PCR_ENTRY_9_8                                                                    (32'h1001a7d0)
`define CLP_PV_REG_PCR_ENTRY_9_9                                                                    (32'h1001a7d4)
`define CLP_PV_REG_PCR_ENTRY_9_10                                                                   (32'h1001a7d8)
`define CLP_PV_REG_PCR_ENTRY_9_11                                                                   (32'h1001a7dc)
`define CLP_PV_REG_PCR_ENTRY_10_0                                                                   (32'h1001a7e0)
`define CLP_PV_REG_PCR_ENTRY_10_1                                                                   (32'h1001a7e4)
`define CLP_PV_REG_PCR_ENTRY_10_2                                                                   (32'h1001a7e8)
`define CLP_PV_REG_PCR_ENTRY_10_3                                                                   (32'h1001a7ec)
`define CLP_PV_REG_PCR_ENTRY_10_4                                                                   (32'h1001a7f0)
`define CLP_PV_REG_PCR_ENTRY_10_5                                                                   (32'h1001a7f4)
`define CLP_PV_REG_PCR_ENTRY_10_6                                                                   (32'h1001a7f8)
`define CLP_PV_REG_PCR_ENTRY_10_7                                                                   (32'h1001a7fc)
`define CLP_PV_REG_PCR_ENTRY_10_8                                                                   (32'h1001a800)
`define CLP_PV_REG_PCR_ENTRY_10_9                                                                   (32'h1001a804)
`define CLP_PV_REG_PCR_ENTRY_10_10                                                                  (32'h1001a808)
`define CLP_PV_REG_PCR_ENTRY_10_11                                                                  (32'h1001a80c)
`define CLP_PV_REG_PCR_ENTRY_11_0                                                                   (32'h1001a810)
`define CLP_PV_REG_PCR_ENTRY_11_1                                                                   (32'h1001a814)
`define CLP_PV_REG_PCR_ENTRY_11_2                                                                   (32'h1001a818)
`define CLP_PV_REG_PCR_ENTRY_11_3                                                                   (32'h1001a81c)
`define CLP_PV_REG_PCR_ENTRY_11_4                                                                   (32'h1001a820)
`define CLP_PV_REG_PCR_ENTRY_11_5                                                                   (32'h1001a824)
`define CLP_PV_REG_PCR_ENTRY_11_6                                                                   (32'h1001a828)
`define CLP_PV_REG_PCR_ENTRY_11_7                                                                   (32'h1001a82c)
`define CLP_PV_REG_PCR_ENTRY_11_8                                                                   (32'h1001a830)
`define CLP_PV_REG_PCR_ENTRY_11_9                                                                   (32'h1001a834)
`define CLP_PV_REG_PCR_ENTRY_11_10                                                                  (32'h1001a838)
`define CLP_PV_REG_PCR_ENTRY_11_11                                                                  (32'h1001a83c)
`define CLP_PV_REG_PCR_ENTRY_12_0                                                                   (32'h1001a840)
`define CLP_PV_REG_PCR_ENTRY_12_1                                                                   (32'h1001a844)
`define CLP_PV_REG_PCR_ENTRY_12_2                                                                   (32'h1001a848)
`define CLP_PV_REG_PCR_ENTRY_12_3                                                                   (32'h1001a84c)
`define CLP_PV_REG_PCR_ENTRY_12_4                                                                   (32'h1001a850)
`define CLP_PV_REG_PCR_ENTRY_12_5                                                                   (32'h1001a854)
`define CLP_PV_REG_PCR_ENTRY_12_6                                                                   (32'h1001a858)
`define CLP_PV_REG_PCR_ENTRY_12_7                                                                   (32'h1001a85c)
`define CLP_PV_REG_PCR_ENTRY_12_8                                                                   (32'h1001a860)
`define CLP_PV_REG_PCR_ENTRY_12_9                                                                   (32'h1001a864)
`define CLP_PV_REG_PCR_ENTRY_12_10                                                                  (32'h1001a868)
`define CLP_PV_REG_PCR_ENTRY_12_11                                                                  (32'h1001a86c)
`define CLP_PV_REG_PCR_ENTRY_13_0                                                                   (32'h1001a870)
`define CLP_PV_REG_PCR_ENTRY_13_1                                                                   (32'h1001a874)
`define CLP_PV_REG_PCR_ENTRY_13_2                                                                   (32'h1001a878)
`define CLP_PV_REG_PCR_ENTRY_13_3                                                                   (32'h1001a87c)
`define CLP_PV_REG_PCR_ENTRY_13_4                                                                   (32'h1001a880)
`define CLP_PV_REG_PCR_ENTRY_13_5                                                                   (32'h1001a884)
`define CLP_PV_REG_PCR_ENTRY_13_6                                                                   (32'h1001a888)
`define CLP_PV_REG_PCR_ENTRY_13_7                                                                   (32'h1001a88c)
`define CLP_PV_REG_PCR_ENTRY_13_8                                                                   (32'h1001a890)
`define CLP_PV_REG_PCR_ENTRY_13_9                                                                   (32'h1001a894)
`define CLP_PV_REG_PCR_ENTRY_13_10                                                                  (32'h1001a898)
`define CLP_PV_REG_PCR_ENTRY_13_11                                                                  (32'h1001a89c)
`define CLP_PV_REG_PCR_ENTRY_14_0                                                                   (32'h1001a8a0)
`define CLP_PV_REG_PCR_ENTRY_14_1                                                                   (32'h1001a8a4)
`define CLP_PV_REG_PCR_ENTRY_14_2                                                                   (32'h1001a8a8)
`define CLP_PV_REG_PCR_ENTRY_14_3                                                                   (32'h1001a8ac)
`define CLP_PV_REG_PCR_ENTRY_14_4                                                                   (32'h1001a8b0)
`define CLP_PV_REG_PCR_ENTRY_14_5                                                                   (32'h1001a8b4)
`define CLP_PV_REG_PCR_ENTRY_14_6                                                                   (32'h1001a8b8)
`define CLP_PV_REG_PCR_ENTRY_14_7                                                                   (32'h1001a8bc)
`define CLP_PV_REG_PCR_ENTRY_14_8                                                                   (32'h1001a8c0)
`define CLP_PV_REG_PCR_ENTRY_14_9                                                                   (32'h1001a8c4)
`define CLP_PV_REG_PCR_ENTRY_14_10                                                                  (32'h1001a8c8)
`define CLP_PV_REG_PCR_ENTRY_14_11                                                                  (32'h1001a8cc)
`define CLP_PV_REG_PCR_ENTRY_15_0                                                                   (32'h1001a8d0)
`define CLP_PV_REG_PCR_ENTRY_15_1                                                                   (32'h1001a8d4)
`define CLP_PV_REG_PCR_ENTRY_15_2                                                                   (32'h1001a8d8)
`define CLP_PV_REG_PCR_ENTRY_15_3                                                                   (32'h1001a8dc)
`define CLP_PV_REG_PCR_ENTRY_15_4                                                                   (32'h1001a8e0)
`define CLP_PV_REG_PCR_ENTRY_15_5                                                                   (32'h1001a8e4)
`define CLP_PV_REG_PCR_ENTRY_15_6                                                                   (32'h1001a8e8)
`define CLP_PV_REG_PCR_ENTRY_15_7                                                                   (32'h1001a8ec)
`define CLP_PV_REG_PCR_ENTRY_15_8                                                                   (32'h1001a8f0)
`define CLP_PV_REG_PCR_ENTRY_15_9                                                                   (32'h1001a8f4)
`define CLP_PV_REG_PCR_ENTRY_15_10                                                                  (32'h1001a8f8)
`define CLP_PV_REG_PCR_ENTRY_15_11                                                                  (32'h1001a8fc)
`define CLP_PV_REG_PCR_ENTRY_16_0                                                                   (32'h1001a900)
`define CLP_PV_REG_PCR_ENTRY_16_1                                                                   (32'h1001a904)
`define CLP_PV_REG_PCR_ENTRY_16_2                                                                   (32'h1001a908)
`define CLP_PV_REG_PCR_ENTRY_16_3                                                                   (32'h1001a90c)
`define CLP_PV_REG_PCR_ENTRY_16_4                                                                   (32'h1001a910)
`define CLP_PV_REG_PCR_ENTRY_16_5                                                                   (32'h1001a914)
`define CLP_PV_REG_PCR_ENTRY_16_6                                                                   (32'h1001a918)
`define CLP_PV_REG_PCR_ENTRY_16_7                                                                   (32'h1001a91c)
`define CLP_PV_REG_PCR_ENTRY_16_8                                                                   (32'h1001a920)
`define CLP_PV_REG_PCR_ENTRY_16_9                                                                   (32'h1001a924)
`define CLP_PV_REG_PCR_ENTRY_16_10                                                                  (32'h1001a928)
`define CLP_PV_REG_PCR_ENTRY_16_11                                                                  (32'h1001a92c)
`define CLP_PV_REG_PCR_ENTRY_17_0                                                                   (32'h1001a930)
`define CLP_PV_REG_PCR_ENTRY_17_1                                                                   (32'h1001a934)
`define CLP_PV_REG_PCR_ENTRY_17_2                                                                   (32'h1001a938)
`define CLP_PV_REG_PCR_ENTRY_17_3                                                                   (32'h1001a93c)
`define CLP_PV_REG_PCR_ENTRY_17_4                                                                   (32'h1001a940)
`define CLP_PV_REG_PCR_ENTRY_17_5                                                                   (32'h1001a944)
`define CLP_PV_REG_PCR_ENTRY_17_6                                                                   (32'h1001a948)
`define CLP_PV_REG_PCR_ENTRY_17_7                                                                   (32'h1001a94c)
`define CLP_PV_REG_PCR_ENTRY_17_8                                                                   (32'h1001a950)
`define CLP_PV_REG_PCR_ENTRY_17_9                                                                   (32'h1001a954)
`define CLP_PV_REG_PCR_ENTRY_17_10                                                                  (32'h1001a958)
`define CLP_PV_REG_PCR_ENTRY_17_11                                                                  (32'h1001a95c)
`define CLP_PV_REG_PCR_ENTRY_18_0                                                                   (32'h1001a960)
`define CLP_PV_REG_PCR_ENTRY_18_1                                                                   (32'h1001a964)
`define CLP_PV_REG_PCR_ENTRY_18_2                                                                   (32'h1001a968)
`define CLP_PV_REG_PCR_ENTRY_18_3                                                                   (32'h1001a96c)
`define CLP_PV_REG_PCR_ENTRY_18_4                                                                   (32'h1001a970)
`define CLP_PV_REG_PCR_ENTRY_18_5                                                                   (32'h1001a974)
`define CLP_PV_REG_PCR_ENTRY_18_6                                                                   (32'h1001a978)
`define CLP_PV_REG_PCR_ENTRY_18_7                                                                   (32'h1001a97c)
`define CLP_PV_REG_PCR_ENTRY_18_8                                                                   (32'h1001a980)
`define CLP_PV_REG_PCR_ENTRY_18_9                                                                   (32'h1001a984)
`define CLP_PV_REG_PCR_ENTRY_18_10                                                                  (32'h1001a988)
`define CLP_PV_REG_PCR_ENTRY_18_11                                                                  (32'h1001a98c)
`define CLP_PV_REG_PCR_ENTRY_19_0                                                                   (32'h1001a990)
`define CLP_PV_REG_PCR_ENTRY_19_1                                                                   (32'h1001a994)
`define CLP_PV_REG_PCR_ENTRY_19_2                                                                   (32'h1001a998)
`define CLP_PV_REG_PCR_ENTRY_19_3                                                                   (32'h1001a99c)
`define CLP_PV_REG_PCR_ENTRY_19_4                                                                   (32'h1001a9a0)
`define CLP_PV_REG_PCR_ENTRY_19_5                                                                   (32'h1001a9a4)
`define CLP_PV_REG_PCR_ENTRY_19_6                                                                   (32'h1001a9a8)
`define CLP_PV_REG_PCR_ENTRY_19_7                                                                   (32'h1001a9ac)
`define CLP_PV_REG_PCR_ENTRY_19_8                                                                   (32'h1001a9b0)
`define CLP_PV_REG_PCR_ENTRY_19_9                                                                   (32'h1001a9b4)
`define CLP_PV_REG_PCR_ENTRY_19_10                                                                  (32'h1001a9b8)
`define CLP_PV_REG_PCR_ENTRY_19_11                                                                  (32'h1001a9bc)
`define CLP_PV_REG_PCR_ENTRY_20_0                                                                   (32'h1001a9c0)
`define CLP_PV_REG_PCR_ENTRY_20_1                                                                   (32'h1001a9c4)
`define CLP_PV_REG_PCR_ENTRY_20_2                                                                   (32'h1001a9c8)
`define CLP_PV_REG_PCR_ENTRY_20_3                                                                   (32'h1001a9cc)
`define CLP_PV_REG_PCR_ENTRY_20_4                                                                   (32'h1001a9d0)
`define CLP_PV_REG_PCR_ENTRY_20_5                                                                   (32'h1001a9d4)
`define CLP_PV_REG_PCR_ENTRY_20_6                                                                   (32'h1001a9d8)
`define CLP_PV_REG_PCR_ENTRY_20_7                                                                   (32'h1001a9dc)
`define CLP_PV_REG_PCR_ENTRY_20_8                                                                   (32'h1001a9e0)
`define CLP_PV_REG_PCR_ENTRY_20_9                                                                   (32'h1001a9e4)
`define CLP_PV_REG_PCR_ENTRY_20_10                                                                  (32'h1001a9e8)
`define CLP_PV_REG_PCR_ENTRY_20_11                                                                  (32'h1001a9ec)
`define CLP_PV_REG_PCR_ENTRY_21_0                                                                   (32'h1001a9f0)
`define CLP_PV_REG_PCR_ENTRY_21_1                                                                   (32'h1001a9f4)
`define CLP_PV_REG_PCR_ENTRY_21_2                                                                   (32'h1001a9f8)
`define CLP_PV_REG_PCR_ENTRY_21_3                                                                   (32'h1001a9fc)
`define CLP_PV_REG_PCR_ENTRY_21_4                                                                   (32'h1001aa00)
`define CLP_PV_REG_PCR_ENTRY_21_5                                                                   (32'h1001aa04)
`define CLP_PV_REG_PCR_ENTRY_21_6                                                                   (32'h1001aa08)
`define CLP_PV_REG_PCR_ENTRY_21_7                                                                   (32'h1001aa0c)
`define CLP_PV_REG_PCR_ENTRY_21_8                                                                   (32'h1001aa10)
`define CLP_PV_REG_PCR_ENTRY_21_9                                                                   (32'h1001aa14)
`define CLP_PV_REG_PCR_ENTRY_21_10                                                                  (32'h1001aa18)
`define CLP_PV_REG_PCR_ENTRY_21_11                                                                  (32'h1001aa1c)
`define CLP_PV_REG_PCR_ENTRY_22_0                                                                   (32'h1001aa20)
`define CLP_PV_REG_PCR_ENTRY_22_1                                                                   (32'h1001aa24)
`define CLP_PV_REG_PCR_ENTRY_22_2                                                                   (32'h1001aa28)
`define CLP_PV_REG_PCR_ENTRY_22_3                                                                   (32'h1001aa2c)
`define CLP_PV_REG_PCR_ENTRY_22_4                                                                   (32'h1001aa30)
`define CLP_PV_REG_PCR_ENTRY_22_5                                                                   (32'h1001aa34)
`define CLP_PV_REG_PCR_ENTRY_22_6                                                                   (32'h1001aa38)
`define CLP_PV_REG_PCR_ENTRY_22_7                                                                   (32'h1001aa3c)
`define CLP_PV_REG_PCR_ENTRY_22_8                                                                   (32'h1001aa40)
`define CLP_PV_REG_PCR_ENTRY_22_9                                                                   (32'h1001aa44)
`define CLP_PV_REG_PCR_ENTRY_22_10                                                                  (32'h1001aa48)
`define CLP_PV_REG_PCR_ENTRY_22_11                                                                  (32'h1001aa4c)
`define CLP_PV_REG_PCR_ENTRY_23_0                                                                   (32'h1001aa50)
`define CLP_PV_REG_PCR_ENTRY_23_1                                                                   (32'h1001aa54)
`define CLP_PV_REG_PCR_ENTRY_23_2                                                                   (32'h1001aa58)
`define CLP_PV_REG_PCR_ENTRY_23_3                                                                   (32'h1001aa5c)
`define CLP_PV_REG_PCR_ENTRY_23_4                                                                   (32'h1001aa60)
`define CLP_PV_REG_PCR_ENTRY_23_5                                                                   (32'h1001aa64)
`define CLP_PV_REG_PCR_ENTRY_23_6                                                                   (32'h1001aa68)
`define CLP_PV_REG_PCR_ENTRY_23_7                                                                   (32'h1001aa6c)
`define CLP_PV_REG_PCR_ENTRY_23_8                                                                   (32'h1001aa70)
`define CLP_PV_REG_PCR_ENTRY_23_9                                                                   (32'h1001aa74)
`define CLP_PV_REG_PCR_ENTRY_23_10                                                                  (32'h1001aa78)
`define CLP_PV_REG_PCR_ENTRY_23_11                                                                  (32'h1001aa7c)
`define CLP_PV_REG_PCR_ENTRY_24_0                                                                   (32'h1001aa80)
`define CLP_PV_REG_PCR_ENTRY_24_1                                                                   (32'h1001aa84)
`define CLP_PV_REG_PCR_ENTRY_24_2                                                                   (32'h1001aa88)
`define CLP_PV_REG_PCR_ENTRY_24_3                                                                   (32'h1001aa8c)
`define CLP_PV_REG_PCR_ENTRY_24_4                                                                   (32'h1001aa90)
`define CLP_PV_REG_PCR_ENTRY_24_5                                                                   (32'h1001aa94)
`define CLP_PV_REG_PCR_ENTRY_24_6                                                                   (32'h1001aa98)
`define CLP_PV_REG_PCR_ENTRY_24_7                                                                   (32'h1001aa9c)
`define CLP_PV_REG_PCR_ENTRY_24_8                                                                   (32'h1001aaa0)
`define CLP_PV_REG_PCR_ENTRY_24_9                                                                   (32'h1001aaa4)
`define CLP_PV_REG_PCR_ENTRY_24_10                                                                  (32'h1001aaa8)
`define CLP_PV_REG_PCR_ENTRY_24_11                                                                  (32'h1001aaac)
`define CLP_PV_REG_PCR_ENTRY_25_0                                                                   (32'h1001aab0)
`define CLP_PV_REG_PCR_ENTRY_25_1                                                                   (32'h1001aab4)
`define CLP_PV_REG_PCR_ENTRY_25_2                                                                   (32'h1001aab8)
`define CLP_PV_REG_PCR_ENTRY_25_3                                                                   (32'h1001aabc)
`define CLP_PV_REG_PCR_ENTRY_25_4                                                                   (32'h1001aac0)
`define CLP_PV_REG_PCR_ENTRY_25_5                                                                   (32'h1001aac4)
`define CLP_PV_REG_PCR_ENTRY_25_6                                                                   (32'h1001aac8)
`define CLP_PV_REG_PCR_ENTRY_25_7                                                                   (32'h1001aacc)
`define CLP_PV_REG_PCR_ENTRY_25_8                                                                   (32'h1001aad0)
`define CLP_PV_REG_PCR_ENTRY_25_9                                                                   (32'h1001aad4)
`define CLP_PV_REG_PCR_ENTRY_25_10                                                                  (32'h1001aad8)
`define CLP_PV_REG_PCR_ENTRY_25_11                                                                  (32'h1001aadc)
`define CLP_PV_REG_PCR_ENTRY_26_0                                                                   (32'h1001aae0)
`define CLP_PV_REG_PCR_ENTRY_26_1                                                                   (32'h1001aae4)
`define CLP_PV_REG_PCR_ENTRY_26_2                                                                   (32'h1001aae8)
`define CLP_PV_REG_PCR_ENTRY_26_3                                                                   (32'h1001aaec)
`define CLP_PV_REG_PCR_ENTRY_26_4                                                                   (32'h1001aaf0)
`define CLP_PV_REG_PCR_ENTRY_26_5                                                                   (32'h1001aaf4)
`define CLP_PV_REG_PCR_ENTRY_26_6                                                                   (32'h1001aaf8)
`define CLP_PV_REG_PCR_ENTRY_26_7                                                                   (32'h1001aafc)
`define CLP_PV_REG_PCR_ENTRY_26_8                                                                   (32'h1001ab00)
`define CLP_PV_REG_PCR_ENTRY_26_9                                                                   (32'h1001ab04)
`define CLP_PV_REG_PCR_ENTRY_26_10                                                                  (32'h1001ab08)
`define CLP_PV_REG_PCR_ENTRY_26_11                                                                  (32'h1001ab0c)
`define CLP_PV_REG_PCR_ENTRY_27_0                                                                   (32'h1001ab10)
`define CLP_PV_REG_PCR_ENTRY_27_1                                                                   (32'h1001ab14)
`define CLP_PV_REG_PCR_ENTRY_27_2                                                                   (32'h1001ab18)
`define CLP_PV_REG_PCR_ENTRY_27_3                                                                   (32'h1001ab1c)
`define CLP_PV_REG_PCR_ENTRY_27_4                                                                   (32'h1001ab20)
`define CLP_PV_REG_PCR_ENTRY_27_5                                                                   (32'h1001ab24)
`define CLP_PV_REG_PCR_ENTRY_27_6                                                                   (32'h1001ab28)
`define CLP_PV_REG_PCR_ENTRY_27_7                                                                   (32'h1001ab2c)
`define CLP_PV_REG_PCR_ENTRY_27_8                                                                   (32'h1001ab30)
`define CLP_PV_REG_PCR_ENTRY_27_9                                                                   (32'h1001ab34)
`define CLP_PV_REG_PCR_ENTRY_27_10                                                                  (32'h1001ab38)
`define CLP_PV_REG_PCR_ENTRY_27_11                                                                  (32'h1001ab3c)
`define CLP_PV_REG_PCR_ENTRY_28_0                                                                   (32'h1001ab40)
`define CLP_PV_REG_PCR_ENTRY_28_1                                                                   (32'h1001ab44)
`define CLP_PV_REG_PCR_ENTRY_28_2                                                                   (32'h1001ab48)
`define CLP_PV_REG_PCR_ENTRY_28_3                                                                   (32'h1001ab4c)
`define CLP_PV_REG_PCR_ENTRY_28_4                                                                   (32'h1001ab50)
`define CLP_PV_REG_PCR_ENTRY_28_5                                                                   (32'h1001ab54)
`define CLP_PV_REG_PCR_ENTRY_28_6                                                                   (32'h1001ab58)
`define CLP_PV_REG_PCR_ENTRY_28_7                                                                   (32'h1001ab5c)
`define CLP_PV_REG_PCR_ENTRY_28_8                                                                   (32'h1001ab60)
`define CLP_PV_REG_PCR_ENTRY_28_9                                                                   (32'h1001ab64)
`define CLP_PV_REG_PCR_ENTRY_28_10                                                                  (32'h1001ab68)
`define CLP_PV_REG_PCR_ENTRY_28_11                                                                  (32'h1001ab6c)
`define CLP_PV_REG_PCR_ENTRY_29_0                                                                   (32'h1001ab70)
`define CLP_PV_REG_PCR_ENTRY_29_1                                                                   (32'h1001ab74)
`define CLP_PV_REG_PCR_ENTRY_29_2                                                                   (32'h1001ab78)
`define CLP_PV_REG_PCR_ENTRY_29_3                                                                   (32'h1001ab7c)
`define CLP_PV_REG_PCR_ENTRY_29_4                                                                   (32'h1001ab80)
`define CLP_PV_REG_PCR_ENTRY_29_5                                                                   (32'h1001ab84)
`define CLP_PV_REG_PCR_ENTRY_29_6                                                                   (32'h1001ab88)
`define CLP_PV_REG_PCR_ENTRY_29_7                                                                   (32'h1001ab8c)
`define CLP_PV_REG_PCR_ENTRY_29_8                                                                   (32'h1001ab90)
`define CLP_PV_REG_PCR_ENTRY_29_9                                                                   (32'h1001ab94)
`define CLP_PV_REG_PCR_ENTRY_29_10                                                                  (32'h1001ab98)
`define CLP_PV_REG_PCR_ENTRY_29_11                                                                  (32'h1001ab9c)
`define CLP_PV_REG_PCR_ENTRY_30_0                                                                   (32'h1001aba0)
`define CLP_PV_REG_PCR_ENTRY_30_1                                                                   (32'h1001aba4)
`define CLP_PV_REG_PCR_ENTRY_30_2                                                                   (32'h1001aba8)
`define CLP_PV_REG_PCR_ENTRY_30_3                                                                   (32'h1001abac)
`define CLP_PV_REG_PCR_ENTRY_30_4                                                                   (32'h1001abb0)
`define CLP_PV_REG_PCR_ENTRY_30_5                                                                   (32'h1001abb4)
`define CLP_PV_REG_PCR_ENTRY_30_6                                                                   (32'h1001abb8)
`define CLP_PV_REG_PCR_ENTRY_30_7                                                                   (32'h1001abbc)
`define CLP_PV_REG_PCR_ENTRY_30_8                                                                   (32'h1001abc0)
`define CLP_PV_REG_PCR_ENTRY_30_9                                                                   (32'h1001abc4)
`define CLP_PV_REG_PCR_ENTRY_30_10                                                                  (32'h1001abc8)
`define CLP_PV_REG_PCR_ENTRY_30_11                                                                  (32'h1001abcc)
`define CLP_PV_REG_PCR_ENTRY_31_0                                                                   (32'h1001abd0)
`define CLP_PV_REG_PCR_ENTRY_31_1                                                                   (32'h1001abd4)
`define CLP_PV_REG_PCR_ENTRY_31_2                                                                   (32'h1001abd8)
`define CLP_PV_REG_PCR_ENTRY_31_3                                                                   (32'h1001abdc)
`define CLP_PV_REG_PCR_ENTRY_31_4                                                                   (32'h1001abe0)
`define CLP_PV_REG_PCR_ENTRY_31_5                                                                   (32'h1001abe4)
`define CLP_PV_REG_PCR_ENTRY_31_6                                                                   (32'h1001abe8)
`define CLP_PV_REG_PCR_ENTRY_31_7                                                                   (32'h1001abec)
`define CLP_PV_REG_PCR_ENTRY_31_8                                                                   (32'h1001abf0)
`define CLP_PV_REG_PCR_ENTRY_31_9                                                                   (32'h1001abf4)
`define CLP_PV_REG_PCR_ENTRY_31_10                                                                  (32'h1001abf8)
`define CLP_PV_REG_PCR_ENTRY_31_11                                                                  (32'h1001abfc)
`define CLP_DV_REG_BASE_ADDR                                                                        (32'h1001c000)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_0                                                            (32'h1001c000)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_1                                                            (32'h1001c004)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_2                                                            (32'h1001c008)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_3                                                            (32'h1001c00c)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_4                                                            (32'h1001c010)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_5                                                            (32'h1001c014)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_6                                                            (32'h1001c018)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_7                                                            (32'h1001c01c)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_8                                                            (32'h1001c020)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_9                                                            (32'h1001c024)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_0                                                      (32'h1001c028)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_1                                                      (32'h1001c02c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_2                                                      (32'h1001c030)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_3                                                      (32'h1001c034)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_4                                                      (32'h1001c038)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_5                                                      (32'h1001c03c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_6                                                      (32'h1001c040)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_7                                                      (32'h1001c044)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_8                                                      (32'h1001c048)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_9                                                      (32'h1001c04c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_10                                                     (32'h1001c050)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_11                                                     (32'h1001c054)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_0                                                      (32'h1001c058)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_1                                                      (32'h1001c05c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_2                                                      (32'h1001c060)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_3                                                      (32'h1001c064)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_4                                                      (32'h1001c068)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_5                                                      (32'h1001c06c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_6                                                      (32'h1001c070)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_7                                                      (32'h1001c074)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_8                                                      (32'h1001c078)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_9                                                      (32'h1001c07c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_10                                                     (32'h1001c080)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_11                                                     (32'h1001c084)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_0                                                      (32'h1001c088)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_1                                                      (32'h1001c08c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_2                                                      (32'h1001c090)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_3                                                      (32'h1001c094)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_4                                                      (32'h1001c098)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_5                                                      (32'h1001c09c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_6                                                      (32'h1001c0a0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_7                                                      (32'h1001c0a4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_8                                                      (32'h1001c0a8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_9                                                      (32'h1001c0ac)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_10                                                     (32'h1001c0b0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_11                                                     (32'h1001c0b4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_0                                                      (32'h1001c0b8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_1                                                      (32'h1001c0bc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_2                                                      (32'h1001c0c0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_3                                                      (32'h1001c0c4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_4                                                      (32'h1001c0c8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_5                                                      (32'h1001c0cc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_6                                                      (32'h1001c0d0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_7                                                      (32'h1001c0d4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_8                                                      (32'h1001c0d8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_9                                                      (32'h1001c0dc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_10                                                     (32'h1001c0e0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_11                                                     (32'h1001c0e4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_0                                                      (32'h1001c0e8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_1                                                      (32'h1001c0ec)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_2                                                      (32'h1001c0f0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_3                                                      (32'h1001c0f4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_4                                                      (32'h1001c0f8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_5                                                      (32'h1001c0fc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_6                                                      (32'h1001c100)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_7                                                      (32'h1001c104)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_8                                                      (32'h1001c108)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_9                                                      (32'h1001c10c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_10                                                     (32'h1001c110)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_11                                                     (32'h1001c114)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_0                                                      (32'h1001c118)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_1                                                      (32'h1001c11c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_2                                                      (32'h1001c120)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_3                                                      (32'h1001c124)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_4                                                      (32'h1001c128)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_5                                                      (32'h1001c12c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_6                                                      (32'h1001c130)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_7                                                      (32'h1001c134)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_8                                                      (32'h1001c138)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_9                                                      (32'h1001c13c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_10                                                     (32'h1001c140)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_11                                                     (32'h1001c144)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_0                                                      (32'h1001c148)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_1                                                      (32'h1001c14c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_2                                                      (32'h1001c150)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_3                                                      (32'h1001c154)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_4                                                      (32'h1001c158)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_5                                                      (32'h1001c15c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_6                                                      (32'h1001c160)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_7                                                      (32'h1001c164)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_8                                                      (32'h1001c168)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_9                                                      (32'h1001c16c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_10                                                     (32'h1001c170)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_11                                                     (32'h1001c174)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_0                                                      (32'h1001c178)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_1                                                      (32'h1001c17c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_2                                                      (32'h1001c180)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_3                                                      (32'h1001c184)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_4                                                      (32'h1001c188)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_5                                                      (32'h1001c18c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_6                                                      (32'h1001c190)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_7                                                      (32'h1001c194)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_8                                                      (32'h1001c198)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_9                                                      (32'h1001c19c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_10                                                     (32'h1001c1a0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_11                                                     (32'h1001c1a4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_0                                                      (32'h1001c1a8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_1                                                      (32'h1001c1ac)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_2                                                      (32'h1001c1b0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_3                                                      (32'h1001c1b4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_4                                                      (32'h1001c1b8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_5                                                      (32'h1001c1bc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_6                                                      (32'h1001c1c0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_7                                                      (32'h1001c1c4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_8                                                      (32'h1001c1c8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_9                                                      (32'h1001c1cc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_10                                                     (32'h1001c1d0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_11                                                     (32'h1001c1d4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_0                                                      (32'h1001c1d8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_1                                                      (32'h1001c1dc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_2                                                      (32'h1001c1e0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_3                                                      (32'h1001c1e4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_4                                                      (32'h1001c1e8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_5                                                      (32'h1001c1ec)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_6                                                      (32'h1001c1f0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_7                                                      (32'h1001c1f4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_8                                                      (32'h1001c1f8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_9                                                      (32'h1001c1fc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_10                                                     (32'h1001c200)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_11                                                     (32'h1001c204)
`define CLP_DV_REG_DATAVAULTCTRL_0                                                                  (32'h1001c208)
`define CLP_DV_REG_DATAVAULTCTRL_1                                                                  (32'h1001c20c)
`define CLP_DV_REG_DATAVAULTCTRL_2                                                                  (32'h1001c210)
`define CLP_DV_REG_DATAVAULTCTRL_3                                                                  (32'h1001c214)
`define CLP_DV_REG_DATAVAULTCTRL_4                                                                  (32'h1001c218)
`define CLP_DV_REG_DATAVAULTCTRL_5                                                                  (32'h1001c21c)
`define CLP_DV_REG_DATAVAULTCTRL_6                                                                  (32'h1001c220)
`define CLP_DV_REG_DATAVAULTCTRL_7                                                                  (32'h1001c224)
`define CLP_DV_REG_DATAVAULTCTRL_8                                                                  (32'h1001c228)
`define CLP_DV_REG_DATAVAULTCTRL_9                                                                  (32'h1001c22c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_0                                                             (32'h1001c230)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_1                                                             (32'h1001c234)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_2                                                             (32'h1001c238)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_3                                                             (32'h1001c23c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_4                                                             (32'h1001c240)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_5                                                             (32'h1001c244)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_6                                                             (32'h1001c248)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_7                                                             (32'h1001c24c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_8                                                             (32'h1001c250)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_9                                                             (32'h1001c254)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_10                                                            (32'h1001c258)
`define CLP_DV_REG_DATA_VAULT_ENTRY_0_11                                                            (32'h1001c25c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_0                                                             (32'h1001c260)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_1                                                             (32'h1001c264)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_2                                                             (32'h1001c268)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_3                                                             (32'h1001c26c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_4                                                             (32'h1001c270)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_5                                                             (32'h1001c274)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_6                                                             (32'h1001c278)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_7                                                             (32'h1001c27c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_8                                                             (32'h1001c280)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_9                                                             (32'h1001c284)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_10                                                            (32'h1001c288)
`define CLP_DV_REG_DATA_VAULT_ENTRY_1_11                                                            (32'h1001c28c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_0                                                             (32'h1001c290)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_1                                                             (32'h1001c294)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_2                                                             (32'h1001c298)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_3                                                             (32'h1001c29c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_4                                                             (32'h1001c2a0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_5                                                             (32'h1001c2a4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_6                                                             (32'h1001c2a8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_7                                                             (32'h1001c2ac)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_8                                                             (32'h1001c2b0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_9                                                             (32'h1001c2b4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_10                                                            (32'h1001c2b8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_2_11                                                            (32'h1001c2bc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_0                                                             (32'h1001c2c0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_1                                                             (32'h1001c2c4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_2                                                             (32'h1001c2c8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_3                                                             (32'h1001c2cc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_4                                                             (32'h1001c2d0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_5                                                             (32'h1001c2d4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_6                                                             (32'h1001c2d8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_7                                                             (32'h1001c2dc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_8                                                             (32'h1001c2e0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_9                                                             (32'h1001c2e4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_10                                                            (32'h1001c2e8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_3_11                                                            (32'h1001c2ec)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_0                                                             (32'h1001c2f0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_1                                                             (32'h1001c2f4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_2                                                             (32'h1001c2f8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_3                                                             (32'h1001c2fc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_4                                                             (32'h1001c300)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_5                                                             (32'h1001c304)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_6                                                             (32'h1001c308)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_7                                                             (32'h1001c30c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_8                                                             (32'h1001c310)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_9                                                             (32'h1001c314)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_10                                                            (32'h1001c318)
`define CLP_DV_REG_DATA_VAULT_ENTRY_4_11                                                            (32'h1001c31c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_0                                                             (32'h1001c320)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_1                                                             (32'h1001c324)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_2                                                             (32'h1001c328)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_3                                                             (32'h1001c32c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_4                                                             (32'h1001c330)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_5                                                             (32'h1001c334)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_6                                                             (32'h1001c338)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_7                                                             (32'h1001c33c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_8                                                             (32'h1001c340)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_9                                                             (32'h1001c344)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_10                                                            (32'h1001c348)
`define CLP_DV_REG_DATA_VAULT_ENTRY_5_11                                                            (32'h1001c34c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_0                                                             (32'h1001c350)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_1                                                             (32'h1001c354)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_2                                                             (32'h1001c358)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_3                                                             (32'h1001c35c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_4                                                             (32'h1001c360)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_5                                                             (32'h1001c364)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_6                                                             (32'h1001c368)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_7                                                             (32'h1001c36c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_8                                                             (32'h1001c370)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_9                                                             (32'h1001c374)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_10                                                            (32'h1001c378)
`define CLP_DV_REG_DATA_VAULT_ENTRY_6_11                                                            (32'h1001c37c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_0                                                             (32'h1001c380)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_1                                                             (32'h1001c384)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_2                                                             (32'h1001c388)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_3                                                             (32'h1001c38c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_4                                                             (32'h1001c390)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_5                                                             (32'h1001c394)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_6                                                             (32'h1001c398)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_7                                                             (32'h1001c39c)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_8                                                             (32'h1001c3a0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_9                                                             (32'h1001c3a4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_10                                                            (32'h1001c3a8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_7_11                                                            (32'h1001c3ac)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_0                                                             (32'h1001c3b0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_1                                                             (32'h1001c3b4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_2                                                             (32'h1001c3b8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_3                                                             (32'h1001c3bc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_4                                                             (32'h1001c3c0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_5                                                             (32'h1001c3c4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_6                                                             (32'h1001c3c8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_7                                                             (32'h1001c3cc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_8                                                             (32'h1001c3d0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_9                                                             (32'h1001c3d4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_10                                                            (32'h1001c3d8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_8_11                                                            (32'h1001c3dc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_0                                                             (32'h1001c3e0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_1                                                             (32'h1001c3e4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_2                                                             (32'h1001c3e8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_3                                                             (32'h1001c3ec)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_4                                                             (32'h1001c3f0)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_5                                                             (32'h1001c3f4)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_6                                                             (32'h1001c3f8)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_7                                                             (32'h1001c3fc)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_8                                                             (32'h1001c400)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_9                                                             (32'h1001c404)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_10                                                            (32'h1001c408)
`define CLP_DV_REG_DATA_VAULT_ENTRY_9_11                                                            (32'h1001c40c)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_0                                                         (32'h1001c410)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_1                                                         (32'h1001c414)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_2                                                         (32'h1001c418)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_3                                                         (32'h1001c41c)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_4                                                         (32'h1001c420)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_5                                                         (32'h1001c424)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_6                                                         (32'h1001c428)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_7                                                         (32'h1001c42c)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_8                                                         (32'h1001c430)
`define CLP_DV_REG_LOCKABLESCRATCHREGCTRL_9                                                         (32'h1001c434)
`define CLP_DV_REG_LOCKABLESCRATCHREG_0                                                             (32'h1001c438)
`define CLP_DV_REG_LOCKABLESCRATCHREG_1                                                             (32'h1001c43c)
`define CLP_DV_REG_LOCKABLESCRATCHREG_2                                                             (32'h1001c440)
`define CLP_DV_REG_LOCKABLESCRATCHREG_3                                                             (32'h1001c444)
`define CLP_DV_REG_LOCKABLESCRATCHREG_4                                                             (32'h1001c448)
`define CLP_DV_REG_LOCKABLESCRATCHREG_5                                                             (32'h1001c44c)
`define CLP_DV_REG_LOCKABLESCRATCHREG_6                                                             (32'h1001c450)
`define CLP_DV_REG_LOCKABLESCRATCHREG_7                                                             (32'h1001c454)
`define CLP_DV_REG_LOCKABLESCRATCHREG_8                                                             (32'h1001c458)
`define CLP_DV_REG_LOCKABLESCRATCHREG_9                                                             (32'h1001c45c)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_0                                                     (32'h1001c460)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_1                                                     (32'h1001c464)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_2                                                     (32'h1001c468)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_3                                                     (32'h1001c46c)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_4                                                     (32'h1001c470)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_5                                                     (32'h1001c474)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_6                                                     (32'h1001c478)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_7                                                     (32'h1001c47c)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0                                                   (32'h1001c480)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1                                                   (32'h1001c484)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2                                                   (32'h1001c488)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3                                                   (32'h1001c48c)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4                                                   (32'h1001c490)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5                                                   (32'h1001c494)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6                                                   (32'h1001c498)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7                                                   (32'h1001c49c)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_0                                                       (32'h1001c4a0)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_1                                                       (32'h1001c4a4)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_2                                                       (32'h1001c4a8)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_3                                                       (32'h1001c4ac)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_4                                                       (32'h1001c4b0)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_5                                                       (32'h1001c4b4)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_6                                                       (32'h1001c4b8)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_7                                                       (32'h1001c4bc)
`define CLP_SHA512_REG_BASE_ADDR                                                                    (32'h10020000)
`define CLP_SHA512_REG_SHA512_NAME_0                                                                (32'h10020000)
`define CLP_SHA512_REG_SHA512_NAME_1                                                                (32'h10020004)
`define CLP_SHA512_REG_SHA512_VERSION_0                                                             (32'h10020008)
`define CLP_SHA512_REG_SHA512_VERSION_1                                                             (32'h1002000c)
`define CLP_SHA512_REG_SHA512_CTRL                                                                  (32'h10020010)
`define CLP_SHA512_REG_SHA512_STATUS                                                                (32'h10020018)
`define CLP_SHA512_REG_SHA512_BLOCK_0                                                               (32'h10020080)
`define CLP_SHA512_REG_SHA512_BLOCK_1                                                               (32'h10020084)
`define CLP_SHA512_REG_SHA512_BLOCK_2                                                               (32'h10020088)
`define CLP_SHA512_REG_SHA512_BLOCK_3                                                               (32'h1002008c)
`define CLP_SHA512_REG_SHA512_BLOCK_4                                                               (32'h10020090)
`define CLP_SHA512_REG_SHA512_BLOCK_5                                                               (32'h10020094)
`define CLP_SHA512_REG_SHA512_BLOCK_6                                                               (32'h10020098)
`define CLP_SHA512_REG_SHA512_BLOCK_7                                                               (32'h1002009c)
`define CLP_SHA512_REG_SHA512_BLOCK_8                                                               (32'h100200a0)
`define CLP_SHA512_REG_SHA512_BLOCK_9                                                               (32'h100200a4)
`define CLP_SHA512_REG_SHA512_BLOCK_10                                                              (32'h100200a8)
`define CLP_SHA512_REG_SHA512_BLOCK_11                                                              (32'h100200ac)
`define CLP_SHA512_REG_SHA512_BLOCK_12                                                              (32'h100200b0)
`define CLP_SHA512_REG_SHA512_BLOCK_13                                                              (32'h100200b4)
`define CLP_SHA512_REG_SHA512_BLOCK_14                                                              (32'h100200b8)
`define CLP_SHA512_REG_SHA512_BLOCK_15                                                              (32'h100200bc)
`define CLP_SHA512_REG_SHA512_BLOCK_16                                                              (32'h100200c0)
`define CLP_SHA512_REG_SHA512_BLOCK_17                                                              (32'h100200c4)
`define CLP_SHA512_REG_SHA512_BLOCK_18                                                              (32'h100200c8)
`define CLP_SHA512_REG_SHA512_BLOCK_19                                                              (32'h100200cc)
`define CLP_SHA512_REG_SHA512_BLOCK_20                                                              (32'h100200d0)
`define CLP_SHA512_REG_SHA512_BLOCK_21                                                              (32'h100200d4)
`define CLP_SHA512_REG_SHA512_BLOCK_22                                                              (32'h100200d8)
`define CLP_SHA512_REG_SHA512_BLOCK_23                                                              (32'h100200dc)
`define CLP_SHA512_REG_SHA512_BLOCK_24                                                              (32'h100200e0)
`define CLP_SHA512_REG_SHA512_BLOCK_25                                                              (32'h100200e4)
`define CLP_SHA512_REG_SHA512_BLOCK_26                                                              (32'h100200e8)
`define CLP_SHA512_REG_SHA512_BLOCK_27                                                              (32'h100200ec)
`define CLP_SHA512_REG_SHA512_BLOCK_28                                                              (32'h100200f0)
`define CLP_SHA512_REG_SHA512_BLOCK_29                                                              (32'h100200f4)
`define CLP_SHA512_REG_SHA512_BLOCK_30                                                              (32'h100200f8)
`define CLP_SHA512_REG_SHA512_BLOCK_31                                                              (32'h100200fc)
`define CLP_SHA512_REG_SHA512_DIGEST_0                                                              (32'h10020100)
`define CLP_SHA512_REG_SHA512_DIGEST_1                                                              (32'h10020104)
`define CLP_SHA512_REG_SHA512_DIGEST_2                                                              (32'h10020108)
`define CLP_SHA512_REG_SHA512_DIGEST_3                                                              (32'h1002010c)
`define CLP_SHA512_REG_SHA512_DIGEST_4                                                              (32'h10020110)
`define CLP_SHA512_REG_SHA512_DIGEST_5                                                              (32'h10020114)
`define CLP_SHA512_REG_SHA512_DIGEST_6                                                              (32'h10020118)
`define CLP_SHA512_REG_SHA512_DIGEST_7                                                              (32'h1002011c)
`define CLP_SHA512_REG_SHA512_DIGEST_8                                                              (32'h10020120)
`define CLP_SHA512_REG_SHA512_DIGEST_9                                                              (32'h10020124)
`define CLP_SHA512_REG_SHA512_DIGEST_10                                                             (32'h10020128)
`define CLP_SHA512_REG_SHA512_DIGEST_11                                                             (32'h1002012c)
`define CLP_SHA512_REG_SHA512_DIGEST_12                                                             (32'h10020130)
`define CLP_SHA512_REG_SHA512_DIGEST_13                                                             (32'h10020134)
`define CLP_SHA512_REG_SHA512_DIGEST_14                                                             (32'h10020138)
`define CLP_SHA512_REG_SHA512_DIGEST_15                                                             (32'h1002013c)
`define CLP_SHA512_REG_SHA512_VAULT_RD_CTRL                                                         (32'h10020600)
`define CLP_SHA512_REG_SHA512_VAULT_RD_STATUS                                                       (32'h10020604)
`define CLP_SHA512_REG_SHA512_KV_WR_CTRL                                                            (32'h10020608)
`define CLP_SHA512_REG_SHA512_KV_WR_STATUS                                                          (32'h1002060c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_0                                                  (32'h10020610)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_1                                                  (32'h10020614)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_2                                                  (32'h10020618)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_3                                                  (32'h1002061c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_4                                                  (32'h10020620)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_5                                                  (32'h10020624)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_6                                                  (32'h10020628)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE_7                                                  (32'h1002062c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_CTRL                                                     (32'h10020630)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_STATUS                                                   (32'h10020634)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_0                                                 (32'h10020638)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_1                                                 (32'h1002063c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_2                                                 (32'h10020640)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_3                                                 (32'h10020644)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_4                                                 (32'h10020648)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_5                                                 (32'h1002064c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_6                                                 (32'h10020650)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_7                                                 (32'h10020654)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_8                                                 (32'h10020658)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_9                                                 (32'h1002065c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_10                                                (32'h10020660)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_11                                                (32'h10020664)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_12                                                (32'h10020668)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_13                                                (32'h1002066c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_14                                                (32'h10020670)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_15                                                (32'h10020674)
`define CLP_SHA512_REG_INTR_BLOCK_RF_START                                                          (32'h10020800)
`define CLP_SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h10020800)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h10020804)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h10020808)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h1002080c)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h10020810)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h10020814)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h10020818)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h1002081c)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h10020820)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h10020900)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h10020904)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h10020908)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h1002090c)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h10020980)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'h10020a00)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'h10020a04)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'h10020a08)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'h10020a0c)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'h10020a10)
`define CLP_SHA256_REG_BASE_ADDR                                                                    (32'h10028000)
`define CLP_SHA256_REG_SHA256_NAME_0                                                                (32'h10028000)
`define CLP_SHA256_REG_SHA256_NAME_1                                                                (32'h10028004)
`define CLP_SHA256_REG_SHA256_VERSION_0                                                             (32'h10028008)
`define CLP_SHA256_REG_SHA256_VERSION_1                                                             (32'h1002800c)
`define CLP_SHA256_REG_SHA256_CTRL                                                                  (32'h10028010)
`define CLP_SHA256_REG_SHA256_STATUS                                                                (32'h10028018)
`define CLP_SHA256_REG_SHA256_BLOCK_0                                                               (32'h10028080)
`define CLP_SHA256_REG_SHA256_BLOCK_1                                                               (32'h10028084)
`define CLP_SHA256_REG_SHA256_BLOCK_2                                                               (32'h10028088)
`define CLP_SHA256_REG_SHA256_BLOCK_3                                                               (32'h1002808c)
`define CLP_SHA256_REG_SHA256_BLOCK_4                                                               (32'h10028090)
`define CLP_SHA256_REG_SHA256_BLOCK_5                                                               (32'h10028094)
`define CLP_SHA256_REG_SHA256_BLOCK_6                                                               (32'h10028098)
`define CLP_SHA256_REG_SHA256_BLOCK_7                                                               (32'h1002809c)
`define CLP_SHA256_REG_SHA256_BLOCK_8                                                               (32'h100280a0)
`define CLP_SHA256_REG_SHA256_BLOCK_9                                                               (32'h100280a4)
`define CLP_SHA256_REG_SHA256_BLOCK_10                                                              (32'h100280a8)
`define CLP_SHA256_REG_SHA256_BLOCK_11                                                              (32'h100280ac)
`define CLP_SHA256_REG_SHA256_BLOCK_12                                                              (32'h100280b0)
`define CLP_SHA256_REG_SHA256_BLOCK_13                                                              (32'h100280b4)
`define CLP_SHA256_REG_SHA256_BLOCK_14                                                              (32'h100280b8)
`define CLP_SHA256_REG_SHA256_BLOCK_15                                                              (32'h100280bc)
`define CLP_SHA256_REG_SHA256_DIGEST_0                                                              (32'h10028100)
`define CLP_SHA256_REG_SHA256_DIGEST_1                                                              (32'h10028104)
`define CLP_SHA256_REG_SHA256_DIGEST_2                                                              (32'h10028108)
`define CLP_SHA256_REG_SHA256_DIGEST_3                                                              (32'h1002810c)
`define CLP_SHA256_REG_SHA256_DIGEST_4                                                              (32'h10028110)
`define CLP_SHA256_REG_SHA256_DIGEST_5                                                              (32'h10028114)
`define CLP_SHA256_REG_SHA256_DIGEST_6                                                              (32'h10028118)
`define CLP_SHA256_REG_SHA256_DIGEST_7                                                              (32'h1002811c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_START                                                          (32'h10028800)
`define CLP_SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h10028800)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h10028804)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h10028808)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h1002880c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h10028810)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h10028814)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h10028818)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h1002881c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h10028820)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h10028900)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h10028904)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h10028908)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h1002890c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h10028980)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'h10028a00)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'h10028a04)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'h10028a08)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'h10028a0c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'h10028a10)
`define CLP_ABR_REG_BASE_ADDR                                                                       (32'h10030000)
`define CLP_ABR_REG_MLDSA_NAME_0                                                                    (32'h10030000)
`define CLP_ABR_REG_MLDSA_NAME_1                                                                    (32'h10030004)
`define CLP_ABR_REG_MLDSA_VERSION_0                                                                 (32'h10030008)
`define CLP_ABR_REG_MLDSA_VERSION_1                                                                 (32'h1003000c)
`define CLP_ABR_REG_MLDSA_CTRL                                                                      (32'h10030010)
`define CLP_ABR_REG_MLDSA_STATUS                                                                    (32'h10030014)
`define CLP_ABR_REG_ABR_ENTROPY_0                                                                   (32'h10030018)
`define CLP_ABR_REG_ABR_ENTROPY_1                                                                   (32'h1003001c)
`define CLP_ABR_REG_ABR_ENTROPY_2                                                                   (32'h10030020)
`define CLP_ABR_REG_ABR_ENTROPY_3                                                                   (32'h10030024)
`define CLP_ABR_REG_ABR_ENTROPY_4                                                                   (32'h10030028)
`define CLP_ABR_REG_ABR_ENTROPY_5                                                                   (32'h1003002c)
`define CLP_ABR_REG_ABR_ENTROPY_6                                                                   (32'h10030030)
`define CLP_ABR_REG_ABR_ENTROPY_7                                                                   (32'h10030034)
`define CLP_ABR_REG_ABR_ENTROPY_8                                                                   (32'h10030038)
`define CLP_ABR_REG_ABR_ENTROPY_9                                                                   (32'h1003003c)
`define CLP_ABR_REG_ABR_ENTROPY_10                                                                  (32'h10030040)
`define CLP_ABR_REG_ABR_ENTROPY_11                                                                  (32'h10030044)
`define CLP_ABR_REG_ABR_ENTROPY_12                                                                  (32'h10030048)
`define CLP_ABR_REG_ABR_ENTROPY_13                                                                  (32'h1003004c)
`define CLP_ABR_REG_ABR_ENTROPY_14                                                                  (32'h10030050)
`define CLP_ABR_REG_ABR_ENTROPY_15                                                                  (32'h10030054)
`define CLP_ABR_REG_MLDSA_SEED_0                                                                    (32'h10030058)
`define CLP_ABR_REG_MLDSA_SEED_1                                                                    (32'h1003005c)
`define CLP_ABR_REG_MLDSA_SEED_2                                                                    (32'h10030060)
`define CLP_ABR_REG_MLDSA_SEED_3                                                                    (32'h10030064)
`define CLP_ABR_REG_MLDSA_SEED_4                                                                    (32'h10030068)
`define CLP_ABR_REG_MLDSA_SEED_5                                                                    (32'h1003006c)
`define CLP_ABR_REG_MLDSA_SEED_6                                                                    (32'h10030070)
`define CLP_ABR_REG_MLDSA_SEED_7                                                                    (32'h10030074)
`define CLP_ABR_REG_MLDSA_SIGN_RND_0                                                                (32'h10030078)
`define CLP_ABR_REG_MLDSA_SIGN_RND_1                                                                (32'h1003007c)
`define CLP_ABR_REG_MLDSA_SIGN_RND_2                                                                (32'h10030080)
`define CLP_ABR_REG_MLDSA_SIGN_RND_3                                                                (32'h10030084)
`define CLP_ABR_REG_MLDSA_SIGN_RND_4                                                                (32'h10030088)
`define CLP_ABR_REG_MLDSA_SIGN_RND_5                                                                (32'h1003008c)
`define CLP_ABR_REG_MLDSA_SIGN_RND_6                                                                (32'h10030090)
`define CLP_ABR_REG_MLDSA_SIGN_RND_7                                                                (32'h10030094)
`define CLP_ABR_REG_MLDSA_MSG_0                                                                     (32'h10030098)
`define CLP_ABR_REG_MLDSA_MSG_1                                                                     (32'h1003009c)
`define CLP_ABR_REG_MLDSA_MSG_2                                                                     (32'h100300a0)
`define CLP_ABR_REG_MLDSA_MSG_3                                                                     (32'h100300a4)
`define CLP_ABR_REG_MLDSA_MSG_4                                                                     (32'h100300a8)
`define CLP_ABR_REG_MLDSA_MSG_5                                                                     (32'h100300ac)
`define CLP_ABR_REG_MLDSA_MSG_6                                                                     (32'h100300b0)
`define CLP_ABR_REG_MLDSA_MSG_7                                                                     (32'h100300b4)
`define CLP_ABR_REG_MLDSA_MSG_8                                                                     (32'h100300b8)
`define CLP_ABR_REG_MLDSA_MSG_9                                                                     (32'h100300bc)
`define CLP_ABR_REG_MLDSA_MSG_10                                                                    (32'h100300c0)
`define CLP_ABR_REG_MLDSA_MSG_11                                                                    (32'h100300c4)
`define CLP_ABR_REG_MLDSA_MSG_12                                                                    (32'h100300c8)
`define CLP_ABR_REG_MLDSA_MSG_13                                                                    (32'h100300cc)
`define CLP_ABR_REG_MLDSA_MSG_14                                                                    (32'h100300d0)
`define CLP_ABR_REG_MLDSA_MSG_15                                                                    (32'h100300d4)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_0                                                              (32'h100300d8)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_1                                                              (32'h100300dc)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_2                                                              (32'h100300e0)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_3                                                              (32'h100300e4)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_4                                                              (32'h100300e8)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_5                                                              (32'h100300ec)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_6                                                              (32'h100300f0)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_7                                                              (32'h100300f4)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_8                                                              (32'h100300f8)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_9                                                              (32'h100300fc)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_10                                                             (32'h10030100)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_11                                                             (32'h10030104)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_12                                                             (32'h10030108)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_13                                                             (32'h1003010c)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_14                                                             (32'h10030110)
`define CLP_ABR_REG_MLDSA_VERIFY_RES_15                                                             (32'h10030114)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_0                                                             (32'h10030118)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_1                                                             (32'h1003011c)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_2                                                             (32'h10030120)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_3                                                             (32'h10030124)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_4                                                             (32'h10030128)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_5                                                             (32'h1003012c)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_6                                                             (32'h10030130)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_7                                                             (32'h10030134)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_8                                                             (32'h10030138)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_9                                                             (32'h1003013c)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_10                                                            (32'h10030140)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_11                                                            (32'h10030144)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_12                                                            (32'h10030148)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_13                                                            (32'h1003014c)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_14                                                            (32'h10030150)
`define CLP_ABR_REG_MLDSA_EXTERNAL_MU_15                                                            (32'h10030154)
`define CLP_ABR_REG_MLDSA_MSG_STROBE                                                                (32'h10030158)
`define CLP_ABR_REG_MLDSA_CTX_CONFIG                                                                (32'h1003015c)
`define CLP_ABR_REG_MLDSA_CTX_0                                                                     (32'h10030160)
`define CLP_ABR_REG_MLDSA_CTX_1                                                                     (32'h10030164)
`define CLP_ABR_REG_MLDSA_CTX_2                                                                     (32'h10030168)
`define CLP_ABR_REG_MLDSA_CTX_3                                                                     (32'h1003016c)
`define CLP_ABR_REG_MLDSA_CTX_4                                                                     (32'h10030170)
`define CLP_ABR_REG_MLDSA_CTX_5                                                                     (32'h10030174)
`define CLP_ABR_REG_MLDSA_CTX_6                                                                     (32'h10030178)
`define CLP_ABR_REG_MLDSA_CTX_7                                                                     (32'h1003017c)
`define CLP_ABR_REG_MLDSA_CTX_8                                                                     (32'h10030180)
`define CLP_ABR_REG_MLDSA_CTX_9                                                                     (32'h10030184)
`define CLP_ABR_REG_MLDSA_CTX_10                                                                    (32'h10030188)
`define CLP_ABR_REG_MLDSA_CTX_11                                                                    (32'h1003018c)
`define CLP_ABR_REG_MLDSA_CTX_12                                                                    (32'h10030190)
`define CLP_ABR_REG_MLDSA_CTX_13                                                                    (32'h10030194)
`define CLP_ABR_REG_MLDSA_CTX_14                                                                    (32'h10030198)
`define CLP_ABR_REG_MLDSA_CTX_15                                                                    (32'h1003019c)
`define CLP_ABR_REG_MLDSA_CTX_16                                                                    (32'h100301a0)
`define CLP_ABR_REG_MLDSA_CTX_17                                                                    (32'h100301a4)
`define CLP_ABR_REG_MLDSA_CTX_18                                                                    (32'h100301a8)
`define CLP_ABR_REG_MLDSA_CTX_19                                                                    (32'h100301ac)
`define CLP_ABR_REG_MLDSA_CTX_20                                                                    (32'h100301b0)
`define CLP_ABR_REG_MLDSA_CTX_21                                                                    (32'h100301b4)
`define CLP_ABR_REG_MLDSA_CTX_22                                                                    (32'h100301b8)
`define CLP_ABR_REG_MLDSA_CTX_23                                                                    (32'h100301bc)
`define CLP_ABR_REG_MLDSA_CTX_24                                                                    (32'h100301c0)
`define CLP_ABR_REG_MLDSA_CTX_25                                                                    (32'h100301c4)
`define CLP_ABR_REG_MLDSA_CTX_26                                                                    (32'h100301c8)
`define CLP_ABR_REG_MLDSA_CTX_27                                                                    (32'h100301cc)
`define CLP_ABR_REG_MLDSA_CTX_28                                                                    (32'h100301d0)
`define CLP_ABR_REG_MLDSA_CTX_29                                                                    (32'h100301d4)
`define CLP_ABR_REG_MLDSA_CTX_30                                                                    (32'h100301d8)
`define CLP_ABR_REG_MLDSA_CTX_31                                                                    (32'h100301dc)
`define CLP_ABR_REG_MLDSA_CTX_32                                                                    (32'h100301e0)
`define CLP_ABR_REG_MLDSA_CTX_33                                                                    (32'h100301e4)
`define CLP_ABR_REG_MLDSA_CTX_34                                                                    (32'h100301e8)
`define CLP_ABR_REG_MLDSA_CTX_35                                                                    (32'h100301ec)
`define CLP_ABR_REG_MLDSA_CTX_36                                                                    (32'h100301f0)
`define CLP_ABR_REG_MLDSA_CTX_37                                                                    (32'h100301f4)
`define CLP_ABR_REG_MLDSA_CTX_38                                                                    (32'h100301f8)
`define CLP_ABR_REG_MLDSA_CTX_39                                                                    (32'h100301fc)
`define CLP_ABR_REG_MLDSA_CTX_40                                                                    (32'h10030200)
`define CLP_ABR_REG_MLDSA_CTX_41                                                                    (32'h10030204)
`define CLP_ABR_REG_MLDSA_CTX_42                                                                    (32'h10030208)
`define CLP_ABR_REG_MLDSA_CTX_43                                                                    (32'h1003020c)
`define CLP_ABR_REG_MLDSA_CTX_44                                                                    (32'h10030210)
`define CLP_ABR_REG_MLDSA_CTX_45                                                                    (32'h10030214)
`define CLP_ABR_REG_MLDSA_CTX_46                                                                    (32'h10030218)
`define CLP_ABR_REG_MLDSA_CTX_47                                                                    (32'h1003021c)
`define CLP_ABR_REG_MLDSA_CTX_48                                                                    (32'h10030220)
`define CLP_ABR_REG_MLDSA_CTX_49                                                                    (32'h10030224)
`define CLP_ABR_REG_MLDSA_CTX_50                                                                    (32'h10030228)
`define CLP_ABR_REG_MLDSA_CTX_51                                                                    (32'h1003022c)
`define CLP_ABR_REG_MLDSA_CTX_52                                                                    (32'h10030230)
`define CLP_ABR_REG_MLDSA_CTX_53                                                                    (32'h10030234)
`define CLP_ABR_REG_MLDSA_CTX_54                                                                    (32'h10030238)
`define CLP_ABR_REG_MLDSA_CTX_55                                                                    (32'h1003023c)
`define CLP_ABR_REG_MLDSA_CTX_56                                                                    (32'h10030240)
`define CLP_ABR_REG_MLDSA_CTX_57                                                                    (32'h10030244)
`define CLP_ABR_REG_MLDSA_CTX_58                                                                    (32'h10030248)
`define CLP_ABR_REG_MLDSA_CTX_59                                                                    (32'h1003024c)
`define CLP_ABR_REG_MLDSA_CTX_60                                                                    (32'h10030250)
`define CLP_ABR_REG_MLDSA_CTX_61                                                                    (32'h10030254)
`define CLP_ABR_REG_MLDSA_CTX_62                                                                    (32'h10030258)
`define CLP_ABR_REG_MLDSA_CTX_63                                                                    (32'h1003025c)
`define CLP_ABR_REG_MLDSA_PUBKEY_BASE_ADDR                                                          (32'h10031000)
`define CLP_ABR_REG_MLDSA_PUBKEY_END_ADDR                                                           (32'h10031a1f)
`define CLP_ABR_REG_MLDSA_SIGNATURE_BASE_ADDR                                                       (32'h10032000)
`define CLP_ABR_REG_MLDSA_SIGNATURE_END_ADDR                                                        (32'h10033213)
`define CLP_ABR_REG_MLDSA_PRIVKEY_OUT_BASE_ADDR                                                     (32'h10034000)
`define CLP_ABR_REG_MLDSA_PRIVKEY_OUT_END_ADDR                                                      (32'h1003531f)
`define CLP_ABR_REG_MLDSA_PRIVKEY_IN_BASE_ADDR                                                      (32'h10036000)
`define CLP_ABR_REG_MLDSA_PRIVKEY_IN_END_ADDR                                                       (32'h1003731f)
`define CLP_ABR_REG_KV_MLDSA_SEED_RD_CTRL                                                           (32'h10038000)
`define CLP_ABR_REG_KV_MLDSA_SEED_RD_STATUS                                                         (32'h10038004)
`define CLP_ABR_REG_INTR_BLOCK_RF_START                                                             (32'h10038100)
`define CLP_ABR_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10038100)
`define CLP_ABR_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10038104)
`define CLP_ABR_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10038108)
`define CLP_ABR_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1003810c)
`define CLP_ABR_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10038110)
`define CLP_ABR_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10038114)
`define CLP_ABR_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10038118)
`define CLP_ABR_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1003811c)
`define CLP_ABR_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10038120)
`define CLP_ABR_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h10038200)
`define CLP_ABR_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10038280)
`define CLP_ABR_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'h10038300)
`define CLP_ABR_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10038304)
`define CLP_ABR_REG_MLKEM_NAME_0                                                                    (32'h10039000)
`define CLP_ABR_REG_MLKEM_NAME_1                                                                    (32'h10039004)
`define CLP_ABR_REG_MLKEM_VERSION_0                                                                 (32'h10039008)
`define CLP_ABR_REG_MLKEM_VERSION_1                                                                 (32'h1003900c)
`define CLP_ABR_REG_MLKEM_CTRL                                                                      (32'h10039010)
`define CLP_ABR_REG_MLKEM_STATUS                                                                    (32'h10039014)
`define CLP_ABR_REG_MLKEM_SEED_D_0                                                                  (32'h10039018)
`define CLP_ABR_REG_MLKEM_SEED_D_1                                                                  (32'h1003901c)
`define CLP_ABR_REG_MLKEM_SEED_D_2                                                                  (32'h10039020)
`define CLP_ABR_REG_MLKEM_SEED_D_3                                                                  (32'h10039024)
`define CLP_ABR_REG_MLKEM_SEED_D_4                                                                  (32'h10039028)
`define CLP_ABR_REG_MLKEM_SEED_D_5                                                                  (32'h1003902c)
`define CLP_ABR_REG_MLKEM_SEED_D_6                                                                  (32'h10039030)
`define CLP_ABR_REG_MLKEM_SEED_D_7                                                                  (32'h10039034)
`define CLP_ABR_REG_MLKEM_SEED_Z_0                                                                  (32'h10039038)
`define CLP_ABR_REG_MLKEM_SEED_Z_1                                                                  (32'h1003903c)
`define CLP_ABR_REG_MLKEM_SEED_Z_2                                                                  (32'h10039040)
`define CLP_ABR_REG_MLKEM_SEED_Z_3                                                                  (32'h10039044)
`define CLP_ABR_REG_MLKEM_SEED_Z_4                                                                  (32'h10039048)
`define CLP_ABR_REG_MLKEM_SEED_Z_5                                                                  (32'h1003904c)
`define CLP_ABR_REG_MLKEM_SEED_Z_6                                                                  (32'h10039050)
`define CLP_ABR_REG_MLKEM_SEED_Z_7                                                                  (32'h10039054)
`define CLP_ABR_REG_MLKEM_SHARED_KEY_0                                                              (32'h10039058)
`define CLP_ABR_REG_MLKEM_SHARED_KEY_1                                                              (32'h1003905c)
`define CLP_ABR_REG_MLKEM_SHARED_KEY_2                                                              (32'h10039060)
`define CLP_ABR_REG_MLKEM_SHARED_KEY_3                                                              (32'h10039064)
`define CLP_ABR_REG_MLKEM_SHARED_KEY_4                                                              (32'h10039068)
`define CLP_ABR_REG_MLKEM_SHARED_KEY_5                                                              (32'h1003906c)
`define CLP_ABR_REG_MLKEM_SHARED_KEY_6                                                              (32'h10039070)
`define CLP_ABR_REG_MLKEM_SHARED_KEY_7                                                              (32'h10039074)
`define CLP_ABR_REG_MLKEM_MSG_BASE_ADDR                                                             (32'h10039080)
`define CLP_ABR_REG_MLKEM_MSG_END_ADDR                                                              (32'h1003909f)
`define CLP_ABR_REG_MLKEM_DECAPS_KEY_BASE_ADDR                                                      (32'h1003a000)
`define CLP_ABR_REG_MLKEM_DECAPS_KEY_END_ADDR                                                       (32'h1003ac5f)
`define CLP_ABR_REG_MLKEM_ENCAPS_KEY_BASE_ADDR                                                      (32'h1003b000)
`define CLP_ABR_REG_MLKEM_ENCAPS_KEY_END_ADDR                                                       (32'h1003b61f)
`define CLP_ABR_REG_MLKEM_CIPHERTEXT_BASE_ADDR                                                      (32'h1003b800)
`define CLP_ABR_REG_MLKEM_CIPHERTEXT_END_ADDR                                                       (32'h1003be1f)
`define CLP_ABR_REG_KV_MLKEM_SEED_RD_CTRL                                                           (32'h1003c000)
`define CLP_ABR_REG_KV_MLKEM_SEED_RD_STATUS                                                         (32'h1003c004)
`define CLP_ABR_REG_KV_MLKEM_MSG_RD_CTRL                                                            (32'h1003c008)
`define CLP_ABR_REG_KV_MLKEM_MSG_RD_STATUS                                                          (32'h1003c00c)
`define CLP_ABR_REG_KV_MLKEM_SHAREDKEY_WR_CTRL                                                      (32'h1003c010)
`define CLP_ABR_REG_KV_MLKEM_SHAREDKEY_WR_STATUS                                                    (32'h1003c014)
`define CLP_KMAC_BASE_ADDR                                                                          (32'h10040000)
`define CLP_KMAC_INTR_STATE                                                                         (32'h10040000)
`define CLP_KMAC_INTR_ENABLE                                                                        (32'h10040004)
`define CLP_KMAC_INTR_TEST                                                                          (32'h10040008)
`define CLP_KMAC_ALERT_TEST                                                                         (32'h1004000c)
`define CLP_KMAC_CFG_REGWEN                                                                         (32'h10040010)
`define CLP_KMAC_CFG_SHADOWED                                                                       (32'h10040014)
`define CLP_KMAC_CMD                                                                                (32'h10040018)
`define CLP_KMAC_STATUS                                                                             (32'h1004001c)
`define CLP_KMAC_PREFIX_0                                                                           (32'h10040020)
`define CLP_KMAC_PREFIX_1                                                                           (32'h10040024)
`define CLP_KMAC_PREFIX_2                                                                           (32'h10040028)
`define CLP_KMAC_PREFIX_3                                                                           (32'h1004002c)
`define CLP_KMAC_PREFIX_4                                                                           (32'h10040030)
`define CLP_KMAC_PREFIX_5                                                                           (32'h10040034)
`define CLP_KMAC_PREFIX_6                                                                           (32'h10040038)
`define CLP_KMAC_PREFIX_7                                                                           (32'h1004003c)
`define CLP_KMAC_PREFIX_8                                                                           (32'h10040040)
`define CLP_KMAC_PREFIX_9                                                                           (32'h10040044)
`define CLP_KMAC_PREFIX_10                                                                          (32'h10040048)
`define CLP_KMAC_ERR_CODE                                                                           (32'h1004004c)
`define CLP_KMAC_STATE_BASE_ADDR                                                                    (32'h10040400)
`define CLP_KMAC_STATE_END_ADDR                                                                     (32'h100404ff)
`define CLP_KMAC_MSG_FIFO_BASE_ADDR                                                                 (32'h10040800)
`define CLP_KMAC_MSG_FIFO_END_ADDR                                                                  (32'h100408ff)
`define CLP_SHA3_BASE_ADDR                                                                          (32'h10041000)
`define CLP_SHA3_SHA3_NAME_0                                                                        (32'h10041000)
`define CLP_SHA3_SHA3_NAME_1                                                                        (32'h10041004)
`define CLP_SHA3_SHA3_VERSION_0                                                                     (32'h10041008)
`define CLP_SHA3_SHA3_VERSION_1                                                                     (32'h1004100c)
`define CLP_SHA3_ALERT_TEST                                                                         (32'h1004101c)
`define CLP_SHA3_CFG_REGWEN                                                                         (32'h10041020)
`define CLP_SHA3_CFG_SHADOWED                                                                       (32'h10041024)
`define CLP_SHA3_CMD                                                                                (32'h10041028)
`define CLP_SHA3_STATUS                                                                             (32'h1004102c)
`define CLP_SHA3_ERR_CODE                                                                           (32'h100410d0)
`define CLP_SHA3_STATE_BASE_ADDR                                                                    (32'h10041200)
`define CLP_SHA3_STATE_END_ADDR                                                                     (32'h100412ff)
`define CLP_SHA3_INTR_BLOCK_RF_START                                                                (32'h10041400)
`define CLP_SHA3_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                     (32'h10041400)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                      (32'h10041404)
`define CLP_SHA3_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                      (32'h10041408)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                  (32'h1004140c)
`define CLP_SHA3_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                  (32'h10041410)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                (32'h10041414)
`define CLP_SHA3_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                (32'h10041418)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                    (32'h1004141c)
`define CLP_SHA3_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                    (32'h10041420)
`define CLP_SHA3_INTR_BLOCK_RF_SHA3_ERROR_INTR_COUNT_R                                              (32'h10041500)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                  (32'h10041504)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                  (32'h10041508)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                  (32'h1004150c)
`define CLP_SHA3_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                          (32'h10041580)
`define CLP_SHA3_INTR_BLOCK_RF_SHA3_ERROR_INTR_COUNT_INCR_R                                         (32'h10041600)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                             (32'h10041604)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                             (32'h10041608)
`define CLP_SHA3_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                             (32'h1004160c)
`define CLP_SHA3_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                     (32'h10041610)
`define CLP_SHA3_MSG_FIFO_BASE_ADDR                                                                 (32'h10041c00)
`define CLP_SHA3_MSG_FIFO_END_ADDR                                                                  (32'h10041cff)
`define CLP_CSRNG_REG_BASE_ADDR                                                                     (32'h20002000)
`define CLP_CSRNG_REG_INTERRUPT_STATE                                                               (32'h20002000)
`define CLP_CSRNG_REG_INTERRUPT_ENABLE                                                              (32'h20002004)
`define CLP_CSRNG_REG_INTERRUPT_TEST                                                                (32'h20002008)
`define CLP_CSRNG_REG_ALERT_TEST                                                                    (32'h2000200c)
`define CLP_CSRNG_REG_REGWEN                                                                        (32'h20002010)
`define CLP_CSRNG_REG_CTRL                                                                          (32'h20002014)
`define CLP_CSRNG_REG_CMD_REQ                                                                       (32'h20002018)
`define CLP_CSRNG_REG_RESEED_INTERVAL                                                               (32'h2000201c)
`define CLP_CSRNG_REG_RESEED_COUNTER_0                                                              (32'h20002020)
`define CLP_CSRNG_REG_RESEED_COUNTER_1                                                              (32'h20002024)
`define CLP_CSRNG_REG_RESEED_COUNTER_2                                                              (32'h20002028)
`define CLP_CSRNG_REG_SW_CMD_STS                                                                    (32'h2000202c)
`define CLP_CSRNG_REG_GENBITS_VLD                                                                   (32'h20002030)
`define CLP_CSRNG_REG_GENBITS                                                                       (32'h20002034)
`define CLP_CSRNG_REG_INT_STATE_READ_ENABLE                                                         (32'h20002038)
`define CLP_CSRNG_REG_INT_STATE_READ_ENABLE_REGWEN                                                  (32'h2000203c)
`define CLP_CSRNG_REG_INT_STATE_NUM                                                                 (32'h20002040)
`define CLP_CSRNG_REG_INT_STATE_VAL                                                                 (32'h20002044)
`define CLP_CSRNG_REG_FIPS_FORCE                                                                    (32'h20002048)
`define CLP_CSRNG_REG_HW_EXC_STS                                                                    (32'h2000204c)
`define CLP_CSRNG_REG_RECOV_ALERT_STS                                                               (32'h20002050)
`define CLP_CSRNG_REG_ERR_CODE                                                                      (32'h20002054)
`define CLP_CSRNG_REG_ERR_CODE_TEST                                                                 (32'h20002058)
`define CLP_CSRNG_REG_MAIN_SM_STATE                                                                 (32'h2000205c)
`define CLP_ENTROPY_SRC_REG_BASE_ADDR                                                               (32'h20003000)
`define CLP_ENTROPY_SRC_REG_INTERRUPT_STATE                                                         (32'h20003000)
`define CLP_ENTROPY_SRC_REG_INTERRUPT_ENABLE                                                        (32'h20003004)
`define CLP_ENTROPY_SRC_REG_INTERRUPT_TEST                                                          (32'h20003008)
`define CLP_ENTROPY_SRC_REG_ALERT_TEST                                                              (32'h2000300c)
`define CLP_ENTROPY_SRC_REG_ME_REGWEN                                                               (32'h20003010)
`define CLP_ENTROPY_SRC_REG_SW_REGUPD                                                               (32'h20003014)
`define CLP_ENTROPY_SRC_REG_REGWEN                                                                  (32'h20003018)
`define CLP_ENTROPY_SRC_REG_REV                                                                     (32'h2000301c)
`define CLP_ENTROPY_SRC_REG_MODULE_ENABLE                                                           (32'h20003020)
`define CLP_ENTROPY_SRC_REG_CONF                                                                    (32'h20003024)
`define CLP_ENTROPY_SRC_REG_ENTROPY_CONTROL                                                         (32'h20003028)
`define CLP_ENTROPY_SRC_REG_ENTROPY_DATA                                                            (32'h2000302c)
`define CLP_ENTROPY_SRC_REG_HEALTH_TEST_WINDOWS                                                     (32'h20003030)
`define CLP_ENTROPY_SRC_REG_REPCNT_THRESHOLDS                                                       (32'h20003034)
`define CLP_ENTROPY_SRC_REG_REPCNTS_THRESHOLDS                                                      (32'h20003038)
`define CLP_ENTROPY_SRC_REG_ADAPTP_HI_THRESHOLDS                                                    (32'h2000303c)
`define CLP_ENTROPY_SRC_REG_ADAPTP_LO_THRESHOLDS                                                    (32'h20003040)
`define CLP_ENTROPY_SRC_REG_BUCKET_THRESHOLDS                                                       (32'h20003044)
`define CLP_ENTROPY_SRC_REG_MARKOV_HI_THRESHOLDS                                                    (32'h20003048)
`define CLP_ENTROPY_SRC_REG_MARKOV_LO_THRESHOLDS                                                    (32'h2000304c)
`define CLP_ENTROPY_SRC_REG_EXTHT_HI_THRESHOLDS                                                     (32'h20003050)
`define CLP_ENTROPY_SRC_REG_EXTHT_LO_THRESHOLDS                                                     (32'h20003054)
`define CLP_ENTROPY_SRC_REG_REPCNT_HI_WATERMARKS                                                    (32'h20003058)
`define CLP_ENTROPY_SRC_REG_REPCNTS_HI_WATERMARKS                                                   (32'h2000305c)
`define CLP_ENTROPY_SRC_REG_ADAPTP_HI_WATERMARKS                                                    (32'h20003060)
`define CLP_ENTROPY_SRC_REG_ADAPTP_LO_WATERMARKS                                                    (32'h20003064)
`define CLP_ENTROPY_SRC_REG_EXTHT_HI_WATERMARKS                                                     (32'h20003068)
`define CLP_ENTROPY_SRC_REG_EXTHT_LO_WATERMARKS                                                     (32'h2000306c)
`define CLP_ENTROPY_SRC_REG_BUCKET_HI_WATERMARKS                                                    (32'h20003070)
`define CLP_ENTROPY_SRC_REG_MARKOV_HI_WATERMARKS                                                    (32'h20003074)
`define CLP_ENTROPY_SRC_REG_MARKOV_LO_WATERMARKS                                                    (32'h20003078)
`define CLP_ENTROPY_SRC_REG_REPCNT_TOTAL_FAILS                                                      (32'h2000307c)
`define CLP_ENTROPY_SRC_REG_REPCNTS_TOTAL_FAILS                                                     (32'h20003080)
`define CLP_ENTROPY_SRC_REG_ADAPTP_HI_TOTAL_FAILS                                                   (32'h20003084)
`define CLP_ENTROPY_SRC_REG_ADAPTP_LO_TOTAL_FAILS                                                   (32'h20003088)
`define CLP_ENTROPY_SRC_REG_BUCKET_TOTAL_FAILS                                                      (32'h2000308c)
`define CLP_ENTROPY_SRC_REG_MARKOV_HI_TOTAL_FAILS                                                   (32'h20003090)
`define CLP_ENTROPY_SRC_REG_MARKOV_LO_TOTAL_FAILS                                                   (32'h20003094)
`define CLP_ENTROPY_SRC_REG_EXTHT_HI_TOTAL_FAILS                                                    (32'h20003098)
`define CLP_ENTROPY_SRC_REG_EXTHT_LO_TOTAL_FAILS                                                    (32'h2000309c)
`define CLP_ENTROPY_SRC_REG_ALERT_THRESHOLD                                                         (32'h200030a0)
`define CLP_ENTROPY_SRC_REG_ALERT_SUMMARY_FAIL_COUNTS                                               (32'h200030a4)
`define CLP_ENTROPY_SRC_REG_ALERT_FAIL_COUNTS                                                       (32'h200030a8)
`define CLP_ENTROPY_SRC_REG_EXTHT_FAIL_COUNTS                                                       (32'h200030ac)
`define CLP_ENTROPY_SRC_REG_FW_OV_CONTROL                                                           (32'h200030b0)
`define CLP_ENTROPY_SRC_REG_FW_OV_SHA3_START                                                        (32'h200030b4)
`define CLP_ENTROPY_SRC_REG_FW_OV_WR_FIFO_FULL                                                      (32'h200030b8)
`define CLP_ENTROPY_SRC_REG_FW_OV_RD_FIFO_OVERFLOW                                                  (32'h200030bc)
`define CLP_ENTROPY_SRC_REG_FW_OV_RD_DATA                                                           (32'h200030c0)
`define CLP_ENTROPY_SRC_REG_FW_OV_WR_DATA                                                           (32'h200030c4)
`define CLP_ENTROPY_SRC_REG_OBSERVE_FIFO_THRESH                                                     (32'h200030c8)
`define CLP_ENTROPY_SRC_REG_OBSERVE_FIFO_DEPTH                                                      (32'h200030cc)
`define CLP_ENTROPY_SRC_REG_DEBUG_STATUS                                                            (32'h200030d0)
`define CLP_ENTROPY_SRC_REG_RECOV_ALERT_STS                                                         (32'h200030d4)
`define CLP_ENTROPY_SRC_REG_ERR_CODE                                                                (32'h200030d8)
`define CLP_ENTROPY_SRC_REG_ERR_CODE_TEST                                                           (32'h200030dc)
`define CLP_ENTROPY_SRC_REG_MAIN_SM_STATE                                                           (32'h200030e0)
`define CLP_MBOX_CSR_BASE_ADDR                                                                      (32'h30020000)
`define CLP_MBOX_CSR_MBOX_LOCK                                                                      (32'h30020000)
`define CLP_MBOX_CSR_MBOX_USER                                                                      (32'h30020004)
`define CLP_MBOX_CSR_MBOX_CMD                                                                       (32'h30020008)
`define CLP_MBOX_CSR_MBOX_DLEN                                                                      (32'h3002000c)
`define CLP_MBOX_CSR_MBOX_DATAIN                                                                    (32'h30020010)
`define CLP_MBOX_CSR_MBOX_DATAOUT                                                                   (32'h30020014)
`define CLP_MBOX_CSR_MBOX_EXECUTE                                                                   (32'h30020018)
`define CLP_MBOX_CSR_MBOX_STATUS                                                                    (32'h3002001c)
`define CLP_MBOX_CSR_MBOX_UNLOCK                                                                    (32'h30020020)
`define CLP_MBOX_CSR_TAP_MODE                                                                       (32'h30020024)
`define CLP_SHA512_ACC_CSR_BASE_ADDR                                                                (32'h30021000)
`define CLP_SHA512_ACC_CSR_LOCK                                                                     (32'h30021000)
`define CLP_SHA512_ACC_CSR_USER                                                                     (32'h30021004)
`define CLP_SHA512_ACC_CSR_MODE                                                                     (32'h30021008)
`define CLP_SHA512_ACC_CSR_START_ADDRESS                                                            (32'h3002100c)
`define CLP_SHA512_ACC_CSR_DLEN                                                                     (32'h30021010)
`define CLP_SHA512_ACC_CSR_DATAIN                                                                   (32'h30021014)
`define CLP_SHA512_ACC_CSR_EXECUTE                                                                  (32'h30021018)
`define CLP_SHA512_ACC_CSR_STATUS                                                                   (32'h3002101c)
`define CLP_SHA512_ACC_CSR_DIGEST_0                                                                 (32'h30021020)
`define CLP_SHA512_ACC_CSR_DIGEST_1                                                                 (32'h30021024)
`define CLP_SHA512_ACC_CSR_DIGEST_2                                                                 (32'h30021028)
`define CLP_SHA512_ACC_CSR_DIGEST_3                                                                 (32'h3002102c)
`define CLP_SHA512_ACC_CSR_DIGEST_4                                                                 (32'h30021030)
`define CLP_SHA512_ACC_CSR_DIGEST_5                                                                 (32'h30021034)
`define CLP_SHA512_ACC_CSR_DIGEST_6                                                                 (32'h30021038)
`define CLP_SHA512_ACC_CSR_DIGEST_7                                                                 (32'h3002103c)
`define CLP_SHA512_ACC_CSR_DIGEST_8                                                                 (32'h30021040)
`define CLP_SHA512_ACC_CSR_DIGEST_9                                                                 (32'h30021044)
`define CLP_SHA512_ACC_CSR_DIGEST_10                                                                (32'h30021048)
`define CLP_SHA512_ACC_CSR_DIGEST_11                                                                (32'h3002104c)
`define CLP_SHA512_ACC_CSR_DIGEST_12                                                                (32'h30021050)
`define CLP_SHA512_ACC_CSR_DIGEST_13                                                                (32'h30021054)
`define CLP_SHA512_ACC_CSR_DIGEST_14                                                                (32'h30021058)
`define CLP_SHA512_ACC_CSR_DIGEST_15                                                                (32'h3002105c)
`define CLP_SHA512_ACC_CSR_CONTROL                                                                  (32'h30021060)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_START                                                      (32'h30021800)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                           (32'h30021800)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R                                            (32'h30021804)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                            (32'h30021808)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                        (32'h3002180c)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                        (32'h30021810)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                      (32'h30021814)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                      (32'h30021818)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                          (32'h3002181c)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                          (32'h30021820)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                        (32'h30021900)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                        (32'h30021904)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                        (32'h30021908)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                        (32'h3002190c)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                (32'h30021980)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                   (32'h30021a00)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                   (32'h30021a04)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                   (32'h30021a08)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                   (32'h30021a0c)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                           (32'h30021a10)
`define CLP_AXI_DMA_REG_BASE_ADDR                                                                   (32'h30022000)
`define CLP_AXI_DMA_REG_ID                                                                          (32'h30022000)
`define CLP_AXI_DMA_REG_CAP                                                                         (32'h30022004)
`define CLP_AXI_DMA_REG_CTRL                                                                        (32'h30022008)
`define CLP_AXI_DMA_REG_STATUS0                                                                     (32'h3002200c)
`define CLP_AXI_DMA_REG_STATUS1                                                                     (32'h30022010)
`define CLP_AXI_DMA_REG_SRC_ADDR_L                                                                  (32'h30022014)
`define CLP_AXI_DMA_REG_SRC_ADDR_H                                                                  (32'h30022018)
`define CLP_AXI_DMA_REG_DST_ADDR_L                                                                  (32'h3002201c)
`define CLP_AXI_DMA_REG_DST_ADDR_H                                                                  (32'h30022020)
`define CLP_AXI_DMA_REG_BYTE_COUNT                                                                  (32'h30022024)
`define CLP_AXI_DMA_REG_BLOCK_SIZE                                                                  (32'h30022028)
`define CLP_AXI_DMA_REG_WRITE_DATA                                                                  (32'h3002202c)
`define CLP_AXI_DMA_REG_READ_DATA                                                                   (32'h30022030)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_START                                                         (32'h30022800)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                              (32'h30022800)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                               (32'h30022804)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                               (32'h30022808)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                           (32'h3002280c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                           (32'h30022810)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                         (32'h30022814)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                         (32'h30022818)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                             (32'h3002281c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                             (32'h30022820)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_CMD_DEC_INTR_COUNT_R                                    (32'h30022900)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_RD_INTR_COUNT_R                                     (32'h30022904)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_WR_INTR_COUNT_R                                     (32'h30022908)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_MBOX_LOCK_INTR_COUNT_R                                  (32'h3002290c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_SHA_LOCK_INTR_COUNT_R                                   (32'h30022910)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_OFLOW_INTR_COUNT_R                                 (32'h30022914)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_UFLOW_INTR_COUNT_R                                 (32'h30022918)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AES_CIF_INTR_COUNT_R                                    (32'h3002291c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_KV_RD_INTR_COUNT_R                                      (32'h30022920)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_KV_RD_LARGE_INTR_COUNT_R                                (32'h30022924)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_TXN_DONE_INTR_COUNT_R                                   (32'h30022980)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_EMPTY_INTR_COUNT_R                                 (32'h30022984)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_EMPTY_INTR_COUNT_R                             (32'h30022988)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_FULL_INTR_COUNT_R                                  (32'h3002298c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_FULL_INTR_COUNT_R                              (32'h30022990)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_CMD_DEC_INTR_COUNT_INCR_R                               (32'h30022a00)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_RD_INTR_COUNT_INCR_R                                (32'h30022a04)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AXI_WR_INTR_COUNT_INCR_R                                (32'h30022a08)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_MBOX_LOCK_INTR_COUNT_INCR_R                             (32'h30022a0c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_SHA_LOCK_INTR_COUNT_INCR_R                              (32'h30022a10)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_OFLOW_INTR_COUNT_INCR_R                            (32'h30022a14)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_FIFO_UFLOW_INTR_COUNT_INCR_R                            (32'h30022a18)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_AES_CIF_INTR_COUNT_INCR_R                               (32'h30022a1c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_KV_RD_INTR_COUNT_INCR_R                                 (32'h30022a20)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_ERROR_KV_RD_LARGE_INTR_COUNT_INCR_R                           (32'h30022a24)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_TXN_DONE_INTR_COUNT_INCR_R                              (32'h30022a28)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_EMPTY_INTR_COUNT_INCR_R                            (32'h30022a2c)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_EMPTY_INTR_COUNT_INCR_R                        (32'h30022a30)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_FULL_INTR_COUNT_INCR_R                             (32'h30022a34)
`define CLP_AXI_DMA_REG_INTR_BLOCK_RF_NOTIF_FIFO_NOT_FULL_INTR_COUNT_INCR_R                         (32'h30022a38)
`define CLP_SOC_IFC_REG_BASE_ADDR                                                                   (32'h30030000)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_FATAL                                                        (32'h30030000)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL                                                    (32'h30030004)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_FATAL                                                        (32'h30030008)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_NON_FATAL                                                    (32'h3003000c)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_ENC                                                          (32'h30030010)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_ENC                                                          (32'h30030014)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                              (32'h30030018)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                              (32'h3003001c)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                              (32'h30030020)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                              (32'h30030024)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                              (32'h30030028)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                              (32'h3003002c)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                              (32'h30030030)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                              (32'h30030034)
`define CLP_SOC_IFC_REG_CPTRA_BOOT_STATUS                                                           (32'h30030038)
`define CLP_SOC_IFC_REG_CPTRA_FLOW_STATUS                                                           (32'h3003003c)
`define CLP_SOC_IFC_REG_CPTRA_RESET_REASON                                                          (32'h30030040)
`define CLP_SOC_IFC_REG_CPTRA_SECURITY_STATE                                                        (32'h30030044)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_0                                                 (32'h30030048)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_1                                                 (32'h3003004c)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_2                                                 (32'h30030050)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_3                                                 (32'h30030054)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_VALID_AXI_USER_4                                                 (32'h30030058)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_0                                                  (32'h3003005c)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_1                                                  (32'h30030060)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_2                                                  (32'h30030064)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_3                                                  (32'h30030068)
`define CLP_SOC_IFC_REG_CPTRA_MBOX_AXI_USER_LOCK_4                                                  (32'h3003006c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_VALID_AXI_USER                                                   (32'h30030070)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_AXI_USER_LOCK                                                    (32'h30030074)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_0                                                           (32'h30030078)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_1                                                           (32'h3003007c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_2                                                           (32'h30030080)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_3                                                           (32'h30030084)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_4                                                           (32'h30030088)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_5                                                           (32'h3003008c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_6                                                           (32'h30030090)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_7                                                           (32'h30030094)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_8                                                           (32'h30030098)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_9                                                           (32'h3003009c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_10                                                          (32'h300300a0)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_11                                                          (32'h300300a4)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_CTRL                                                             (32'h300300a8)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_STATUS                                                           (32'h300300ac)
`define CLP_SOC_IFC_REG_CPTRA_FUSE_WR_DONE                                                          (32'h300300b0)
`define CLP_SOC_IFC_REG_CPTRA_TIMER_CONFIG                                                          (32'h300300b4)
`define CLP_SOC_IFC_REG_CPTRA_BOOTFSM_GO                                                            (32'h300300b8)
`define CLP_SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG                                                 (32'h300300bc)
`define CLP_SOC_IFC_REG_CPTRA_CLK_GATING_EN                                                         (32'h300300c0)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_0                                                 (32'h300300c4)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_1                                                 (32'h300300c8)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                                (32'h300300cc)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                                (32'h300300d0)
`define CLP_SOC_IFC_REG_CPTRA_HW_REV_ID                                                             (32'h300300d4)
`define CLP_SOC_IFC_REG_CPTRA_FW_REV_ID_0                                                           (32'h300300d8)
`define CLP_SOC_IFC_REG_CPTRA_FW_REV_ID_1                                                           (32'h300300dc)
`define CLP_SOC_IFC_REG_CPTRA_HW_CONFIG                                                             (32'h300300e0)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER1_EN                                                         (32'h300300e4)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER1_CTRL                                                       (32'h300300e8)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_0                                           (32'h300300ec)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER1_TIMEOUT_PERIOD_1                                           (32'h300300f0)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER2_EN                                                         (32'h300300f4)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER2_CTRL                                                       (32'h300300f8)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_0                                           (32'h300300fc)
`define CLP_SOC_IFC_REG_CPTRA_WDT_TIMER2_TIMEOUT_PERIOD_1                                           (32'h30030100)
`define CLP_SOC_IFC_REG_CPTRA_WDT_STATUS                                                            (32'h30030104)
`define CLP_SOC_IFC_REG_CPTRA_FUSE_VALID_AXI_USER                                                   (32'h30030108)
`define CLP_SOC_IFC_REG_CPTRA_FUSE_AXI_USER_LOCK                                                    (32'h3003010c)
`define CLP_SOC_IFC_REG_CPTRA_WDT_CFG_0                                                             (32'h30030110)
`define CLP_SOC_IFC_REG_CPTRA_WDT_CFG_1                                                             (32'h30030114)
`define CLP_SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0                                                (32'h30030118)
`define CLP_SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1                                                (32'h3003011c)
`define CLP_SOC_IFC_REG_CPTRA_RSVD_REG_0                                                            (32'h30030120)
`define CLP_SOC_IFC_REG_CPTRA_RSVD_REG_1                                                            (32'h30030124)
`define CLP_SOC_IFC_REG_CPTRA_HW_CAPABILITIES                                                       (32'h30030128)
`define CLP_SOC_IFC_REG_CPTRA_FW_CAPABILITIES                                                       (32'h3003012c)
`define CLP_SOC_IFC_REG_CPTRA_CAP_LOCK                                                              (32'h30030130)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_0                                                       (32'h30030140)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_1                                                       (32'h30030144)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_2                                                       (32'h30030148)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_3                                                       (32'h3003014c)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_4                                                       (32'h30030150)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_5                                                       (32'h30030154)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_6                                                       (32'h30030158)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_7                                                       (32'h3003015c)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_8                                                       (32'h30030160)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_9                                                       (32'h30030164)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_10                                                      (32'h30030168)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_11                                                      (32'h3003016c)
`define CLP_SOC_IFC_REG_CPTRA_OWNER_PK_HASH_LOCK                                                    (32'h30030170)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_0                                                             (32'h30030200)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_1                                                             (32'h30030204)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_2                                                             (32'h30030208)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_3                                                             (32'h3003020c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_4                                                             (32'h30030210)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_5                                                             (32'h30030214)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_6                                                             (32'h30030218)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_7                                                             (32'h3003021c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_8                                                             (32'h30030220)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_9                                                             (32'h30030224)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_10                                                            (32'h30030228)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_11                                                            (32'h3003022c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_12                                                            (32'h30030230)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_13                                                            (32'h30030234)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_14                                                            (32'h30030238)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_15                                                            (32'h3003023c)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_0                                                        (32'h30030240)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_1                                                        (32'h30030244)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_2                                                        (32'h30030248)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_3                                                        (32'h3003024c)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_4                                                        (32'h30030250)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_5                                                        (32'h30030254)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_6                                                        (32'h30030258)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_7                                                        (32'h3003025c)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_0                                                       (32'h30030260)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_1                                                       (32'h30030264)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_2                                                       (32'h30030268)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_3                                                       (32'h3003026c)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_4                                                       (32'h30030270)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_5                                                       (32'h30030274)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_6                                                       (32'h30030278)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_7                                                       (32'h3003027c)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_8                                                       (32'h30030280)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_9                                                       (32'h30030284)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_10                                                      (32'h30030288)
`define CLP_SOC_IFC_REG_FUSE_VENDOR_PK_HASH_11                                                      (32'h3003028c)
`define CLP_SOC_IFC_REG_FUSE_ECC_REVOCATION                                                         (32'h30030290)
`define CLP_SOC_IFC_REG_FUSE_FMC_KEY_MANIFEST_SVN                                                   (32'h300302b4)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_0                                                          (32'h300302b8)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_1                                                          (32'h300302bc)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_2                                                          (32'h300302c0)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_3                                                          (32'h300302c4)
`define CLP_SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE                                                  (32'h300302c8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_0                                                     (32'h300302cc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_1                                                     (32'h300302d0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_2                                                     (32'h300302d4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_3                                                     (32'h300302d8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_4                                                     (32'h300302dc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_5                                                     (32'h300302e0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6                                                     (32'h300302e4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7                                                     (32'h300302e8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8                                                     (32'h300302ec)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9                                                     (32'h300302f0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10                                                    (32'h300302f4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_11                                                    (32'h300302f8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_12                                                    (32'h300302fc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_13                                                    (32'h30030300)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_14                                                    (32'h30030304)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_15                                                    (32'h30030308)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_16                                                    (32'h3003030c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_17                                                    (32'h30030310)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_18                                                    (32'h30030314)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_19                                                    (32'h30030318)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_20                                                    (32'h3003031c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_21                                                    (32'h30030320)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_22                                                    (32'h30030324)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_23                                                    (32'h30030328)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                                  (32'h3003032c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                                  (32'h30030330)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                                  (32'h30030334)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                                  (32'h30030338)
`define CLP_SOC_IFC_REG_FUSE_LMS_REVOCATION                                                         (32'h30030340)
`define CLP_SOC_IFC_REG_FUSE_MLDSA_REVOCATION                                                       (32'h30030344)
`define CLP_SOC_IFC_REG_FUSE_SOC_STEPPING_ID                                                        (32'h30030348)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_0                                               (32'h3003034c)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_1                                               (32'h30030350)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_2                                               (32'h30030354)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_3                                               (32'h30030358)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_4                                               (32'h3003035c)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_5                                               (32'h30030360)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_6                                               (32'h30030364)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_7                                               (32'h30030368)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_8                                               (32'h3003036c)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_9                                               (32'h30030370)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_10                                              (32'h30030374)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_11                                              (32'h30030378)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_12                                              (32'h3003037c)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_13                                              (32'h30030380)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_14                                              (32'h30030384)
`define CLP_SOC_IFC_REG_FUSE_MANUF_DBG_UNLOCK_TOKEN_15                                              (32'h30030388)
`define CLP_SOC_IFC_REG_FUSE_PQC_KEY_TYPE                                                           (32'h3003038c)
`define CLP_SOC_IFC_REG_FUSE_SOC_MANIFEST_SVN_0                                                     (32'h30030390)
`define CLP_SOC_IFC_REG_FUSE_SOC_MANIFEST_SVN_1                                                     (32'h30030394)
`define CLP_SOC_IFC_REG_FUSE_SOC_MANIFEST_SVN_2                                                     (32'h30030398)
`define CLP_SOC_IFC_REG_FUSE_SOC_MANIFEST_SVN_3                                                     (32'h3003039c)
`define CLP_SOC_IFC_REG_FUSE_SOC_MANIFEST_MAX_SVN                                                   (32'h300303a0)
`define CLP_SOC_IFC_REG_FUSE_HEK_SEED_0                                                             (32'h300303c0)
`define CLP_SOC_IFC_REG_FUSE_HEK_SEED_1                                                             (32'h300303c4)
`define CLP_SOC_IFC_REG_FUSE_HEK_SEED_2                                                             (32'h300303c8)
`define CLP_SOC_IFC_REG_FUSE_HEK_SEED_3                                                             (32'h300303cc)
`define CLP_SOC_IFC_REG_FUSE_HEK_SEED_4                                                             (32'h300303d0)
`define CLP_SOC_IFC_REG_FUSE_HEK_SEED_5                                                             (32'h300303d4)
`define CLP_SOC_IFC_REG_FUSE_HEK_SEED_6                                                             (32'h300303d8)
`define CLP_SOC_IFC_REG_FUSE_HEK_SEED_7                                                             (32'h300303dc)
`define CLP_SOC_IFC_REG_SS_CALIPTRA_BASE_ADDR_L                                                     (32'h30030500)
`define CLP_SOC_IFC_REG_SS_CALIPTRA_BASE_ADDR_H                                                     (32'h30030504)
`define CLP_SOC_IFC_REG_SS_MCI_BASE_ADDR_L                                                          (32'h30030508)
`define CLP_SOC_IFC_REG_SS_MCI_BASE_ADDR_H                                                          (32'h3003050c)
`define CLP_SOC_IFC_REG_SS_RECOVERY_IFC_BASE_ADDR_L                                                 (32'h30030510)
`define CLP_SOC_IFC_REG_SS_RECOVERY_IFC_BASE_ADDR_H                                                 (32'h30030514)
`define CLP_SOC_IFC_REG_SS_OTP_FC_BASE_ADDR_L                                                       (32'h30030518)
`define CLP_SOC_IFC_REG_SS_OTP_FC_BASE_ADDR_H                                                       (32'h3003051c)
`define CLP_SOC_IFC_REG_SS_UDS_SEED_BASE_ADDR_L                                                     (32'h30030520)
`define CLP_SOC_IFC_REG_SS_UDS_SEED_BASE_ADDR_H                                                     (32'h30030524)
`define CLP_SOC_IFC_REG_SS_PROD_DEBUG_UNLOCK_AUTH_PK_HASH_REG_BANK_OFFSET                           (32'h30030528)
`define CLP_SOC_IFC_REG_SS_NUM_OF_PROD_DEBUG_UNLOCK_AUTH_PK_HASHES                                  (32'h3003052c)
`define CLP_SOC_IFC_REG_SS_DEBUG_INTENT                                                             (32'h30030530)
`define CLP_SOC_IFC_REG_SS_CALIPTRA_DMA_AXI_USER                                                    (32'h30030534)
`define CLP_SOC_IFC_REG_SS_EXTERNAL_STAGING_AREA_BASE_ADDR_L                                        (32'h30030538)
`define CLP_SOC_IFC_REG_SS_EXTERNAL_STAGING_AREA_BASE_ADDR_H                                        (32'h3003053c)
`define CLP_SOC_IFC_REG_SS_KEY_RELEASE_BASE_ADDR_L                                                  (32'h30030540)
`define CLP_SOC_IFC_REG_SS_KEY_RELEASE_BASE_ADDR_H                                                  (32'h30030544)
`define CLP_SOC_IFC_REG_SS_KEY_RELEASE_SIZE                                                         (32'h30030548)
`define CLP_SOC_IFC_REG_SS_OCP_LOCK_CTRL                                                            (32'h3003054c)
`define CLP_SOC_IFC_REG_SS_STRAP_GENERIC_0                                                          (32'h300305a0)
`define CLP_SOC_IFC_REG_SS_STRAP_GENERIC_1                                                          (32'h300305a4)
`define CLP_SOC_IFC_REG_SS_STRAP_GENERIC_2                                                          (32'h300305a8)
`define CLP_SOC_IFC_REG_SS_STRAP_GENERIC_3                                                          (32'h300305ac)
`define CLP_SOC_IFC_REG_SS_DBG_SERVICE_REG_REQ                                                      (32'h300305c0)
`define CLP_SOC_IFC_REG_SS_DBG_SERVICE_REG_RSP                                                      (32'h300305c4)
`define CLP_SOC_IFC_REG_SS_SOC_DBG_UNLOCK_LEVEL_0                                                   (32'h300305c8)
`define CLP_SOC_IFC_REG_SS_SOC_DBG_UNLOCK_LEVEL_1                                                   (32'h300305cc)
`define CLP_SOC_IFC_REG_SS_GENERIC_FW_EXEC_CTRL_0                                                   (32'h300305d0)
`define CLP_SOC_IFC_REG_SS_GENERIC_FW_EXEC_CTRL_1                                                   (32'h300305d4)
`define CLP_SOC_IFC_REG_SS_GENERIC_FW_EXEC_CTRL_2                                                   (32'h300305d8)
`define CLP_SOC_IFC_REG_SS_GENERIC_FW_EXEC_CTRL_3                                                   (32'h300305dc)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_0                                                          (32'h30030600)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_1                                                          (32'h30030604)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_2                                                          (32'h30030608)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_3                                                          (32'h3003060c)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_4                                                          (32'h30030610)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_5                                                          (32'h30030614)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_6                                                          (32'h30030618)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_7                                                          (32'h3003061c)
`define CLP_SOC_IFC_REG_INTERNAL_ICCM_LOCK                                                          (32'h30030620)
`define CLP_SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET                                                    (32'h30030624)
`define CLP_SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES                                        (32'h30030628)
`define CLP_SOC_IFC_REG_INTERNAL_NMI_VECTOR                                                         (32'h3003062c)
`define CLP_SOC_IFC_REG_INTERNAL_HW_ERROR_FATAL_MASK                                                (32'h30030630)
`define CLP_SOC_IFC_REG_INTERNAL_HW_ERROR_NON_FATAL_MASK                                            (32'h30030634)
`define CLP_SOC_IFC_REG_INTERNAL_FW_ERROR_FATAL_MASK                                                (32'h30030638)
`define CLP_SOC_IFC_REG_INTERNAL_FW_ERROR_NON_FATAL_MASK                                            (32'h3003063c)
`define CLP_SOC_IFC_REG_INTERNAL_RV_MTIME_L                                                         (32'h30030640)
`define CLP_SOC_IFC_REG_INTERNAL_RV_MTIME_H                                                         (32'h30030644)
`define CLP_SOC_IFC_REG_INTERNAL_RV_MTIMECMP_L                                                      (32'h30030648)
`define CLP_SOC_IFC_REG_INTERNAL_RV_MTIMECMP_H                                                      (32'h3003064c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_START                                                         (32'h30030800)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                              (32'h30030800)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                               (32'h30030804)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                               (32'h30030808)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                           (32'h3003080c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                           (32'h30030810)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                         (32'h30030814)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                         (32'h30030818)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                             (32'h3003081c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                             (32'h30030820)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                   (32'h30030900)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_R                                    (32'h30030904)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_R                                   (32'h30030908)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_R                                   (32'h3003090c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_R                               (32'h30030910)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_R                               (32'h30030914)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_R                         (32'h30030918)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_R                         (32'h3003091c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_R                                  (32'h30030980)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_R                               (32'h30030984)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                               (32'h30030988)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_R                                  (32'h3003098c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SOC_REQ_LOCK_INTR_COUNT_R                               (32'h30030990)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_R                              (32'h30030994)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                              (32'h30030a00)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R                               (32'h30030a04)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R                              (32'h30030a08)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R                              (32'h30030a0c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R                          (32'h30030a10)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R                          (32'h30030a14)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER1_TIMEOUT_INTR_COUNT_INCR_R                    (32'h30030a18)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_WDT_TIMER2_TIMEOUT_INTR_COUNT_INCR_R                    (32'h30030a1c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R                             (32'h30030a20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R                          (32'h30030a24)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                          (32'h30030a28)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SCAN_MODE_INTR_COUNT_INCR_R                             (32'h30030a2c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_SOC_REQ_LOCK_INTR_COUNT_INCR_R                          (32'h30030a30)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GEN_IN_TOGGLE_INTR_COUNT_INCR_R                         (32'h30030a34)
`define CLP_MBOX_SRAM_BASE_ADDR                                                                     (32'h30040000)
`define CLP_MBOX_SRAM_END_ADDR                                                                      (32'h30043fff)


`endif