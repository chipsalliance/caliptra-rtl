// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//

`include "caliptra_prim_assert.sv";

module axi_adapter_sram
    import axi_pkg::*;
    import caliptra_prim_mubi_pkg::mubi4_t;
#(
    parameter int SramAw            = 12,
    parameter int SramDw            = 32, // Must be multiple of the TL width
    parameter int Outstanding       = 1,  // Only one request is accepted
    parameter bit ByteAccess        = 1,  // 1: Enables sub-word write transactions. Note that this
                                            //    results in read-modify-write operations for integrity
                                            //    re-generation if EnableDataIntgPt is set to 1.
    parameter bit ErrOnWrite        = 0,  // 1: Writelogic           win_dv,
    logic [AW-1:0]  win_addr,
    logic           win_write,
    //logic [UW-1:0]  win_user,
    logic [IW-1:0]  win_id,
    logic [DW-1:0]  win_wdata,
    logic [BC-1:0]  win_wstrb,
    logic [DW-1:0]  win_rdata,
    logic           win_last,
    logic           win_hld,
    logic           win_err,s not allowed, automatically error
    parameter bit ErrOnRead         = 0,  // 1: Reads not allowed, automatically error
    //parameter bit CmdIntgCheck      = 0,  // 1: Enable command integrity check
    //parameter bit EnableRspIntgGen  = 0,  // 1: Generate response integrity
    //parameter bit EnableDataIntgGen = 0,  // 1: Generate response data integrity
    //parameter bit EnableDataIntgPt  = 0,  // 1: Passthrough command/response data integrity
    //parameter bit SecFifoPtr        = 0,  // 1: Duplicated fifo pointers
    localparam int WidthMult        = SramDw / axi_pkg::AXI_DW,
    //localparam int IntgWidth        = tlul_pkg::DataIntgWidth * WidthMult,
    //localparam int DataOutW         = EnableDataIntgPt ? SramDw + IntgWidth : SramDw
    localparam int DataOutW         = SramDw;
) (
    input clk_i, 
    input rst_ni,

    // AXI interface
    input  logic                        axi_dv,
    input  logic [axi_pkg::AXI_AW-1:0]  axi_addr,
    input  logic                        axi_write,
    input  logic [axi_pkg::AXI_IW-1:0]  axi_id,
    input  logic [axi_pkg::AXI_DW-1:0]  axi_wdata,
    input  logic [axi_pkg::AXI_BC-1:0]  axi_wstrb,
    output logic [axi_pkg::AXI_DW-1:0]  axi_rdata,
    input  logic                        axi_last,
    output logic                        axi_hld,
    output logic                        axi_err,

    // Control interface
    input  mubi4_t                      en_ifetch_i,

    // SRAM interface
    output logic                        req_o,
    output mubi4_t                      req_type_o,
    input                               gnt_i,
    output logic                        we_o,
    output logic [SramAw-1:0]           addr_o,
    output logic [DataOutW-1:0]         wdata_o,
    output logic [DataOutW-1:0]         wmask_o,
    //output logic                        intg_error_o,
    input        [DataOutW-1:0]         rdata_i,
    input                               rvalid_i,
    input        [1:0]                  rerror_i, // 2 bit error [1]: Uncorrectable, [0]: Correctable
    output logic                        rmw_in_progress_o
);

    localparam int SramByte = SramDw/8;
    localparam int DataBitWidth = caliptra_prim_util_pkg::vbits(SramByte);
    localparam int WoffsetWidth = (SramByte == axi_pkg::AXI_BC) ? 1 :
                                    DataBitWidth - caliptra_prim_util_pkg::vbits(axi_pkg::AXI_BC);

    logic error_det; // Internal protocol error checker
    logic error_internal; // Internal protocol error checker
    logic wr_attr_error;
    //logic instr_error; //TODO
    logic wr_vld_error;
    logic rd_vld_error;
    logic rsp_fifo_error;
    //logic intg_error;
    logic axi_error;

    // wr_attr_error: Check if the request size, strb are permitted.
    //    Basic check of size, mask, addr align is done in tlul_err module.
    //    Here it checks any partial write if ByteAccess isn't allowed.
    assign wr_attr_error = (axi_write) ? ((ByteAccess == 0) ? (axi_wstrb != '1) : 1'b0) : 1'b0;

    // TODO: how does this apply to AXI -- instruction type?
    /*
    // An instruction type transaction is only valid if en_ifetch is enabled
    // If the instruction type is completely invalid, also considered an instruction error
    assign instr_error = prim_mubi_pkg::mubi4_test_invalid(tl_i.a_user.instr_type) |
    (prim_mubi_pkg::mubi4_test_true_strict(tl_i.a_user.instr_type) &
    prim_mubi_pkg::mubi4_test_false_loose(en_ifetch_i));
     */                             

    if (ErrOnWrite == 1) begin : gen_no_writes
       assign wr_vld_error = axi_write != 1'b0;
    end else begin : gen_writes_allowed
       assign wr_vld_error = 1'b0;
    end
    
    if (ErrOnRead == 1) begin: gen_no_reads
       assign rd_vld_error = core_write == 1'b0;
    end else begin : gen_reads_allowed
       assign rd_vld_error = 1'b0;
    end

    //TODO: equiv of tlul_protocol check
    // COpyinge existing tlul code for now
    // tlul protocol check
    tlul_err u_err (
        .clk_i,
        .rst_ni,
        .tl_i(tl_i),
        .err_o (tlul_error)
    );

    // error return is transactional and thus does not used the "latched" intg_err signal
    assign error_det = wr_attr_error | wr_vld_error | rd_vld_error | //instr_error |
                            tlul_error;//    | intg_error;

    typedef struct packed {
        logic [axi_pkg::AXI_BC-1:0] wstrb ; // Byte mask within the AXI word
        logic [WoffsetWidth-1:0]    woffset ; // Offset of the TL-UL word within the SRAM word
    } sram_req_t ;

    typedef struct packed {
        logic                       write;
        logic [axi_pkg::AXI_BC-1:0] wstrb;
        logic [axi_pkg::AXI_IW-1:0] id;
        logic                       error;
    } req_t;

    typedef struct packed {
        logic [axi_pkg::AXI_DW-1:0] data;
        logic                       error; 
    } rsp_t;
                            
    localparam int SramReqFifoWidth = $bits(sram_req_t) ;
    localparam int ReqFifoWidth = $bits(req_t) ;
    localparam int RspFifoWidth = $bits(rsp_t) ;

    // FIFO signal in case OutStand is greater than 1
    // If request is latched, {write, source} is pushed to req fifo.
    // Req fifo is popped when axi_dv is asserted and axi_hld is 0.
    // axi_vld is asserted if it is write request or rsp fifo not empty if read.
    logic reqfifo_wvalid, reqfifo_wready;
    logic reqfifo_rvalid, reqfifo_rready;
    req_t reqfifo_wdata,  reqfifo_rdata;

    logic sramreqfifo_wvalid, sramreqfifo_wready;
    logic sramreqfifo_rready;
    sram_req_t sramreqfifo_wdata, sramreqfifo_rdata;

    logic rspfifo_wvalid, rspfifo_wready;
    logic rspfifo_rvalid, rspfifo_rready;
    rsp_t rspfifo_wdata,  rspfifo_rdata;

    logic a_ack, d_ack, sram_ack;
    assign a_ack    = axi_dv & ~axi_hld;
    assign d_ack    = axi_dv & ~ axi_hld;
    assign sram_ack = req_o & gnt_i;

    // Valid handling
    logic d_valid, d_error;
    always_comb begin
        d_valid = 1'b0;
        if (reqfifo_rvalid) begin
            if (reqfifo_rdata.error) begin
                // Return error response. Assume no request went out to SRAM
                d_valid = 1'b1;
            end else if (!reqfifo_rdata.write) begin // Read
                d_valid = rspfifo_rvalid;
            end else begin
                // Write without error
                d_valid = 1'b1;
            end
        end else begin
            d_valid = 1'b0;
        end
    end

    always_comb begin
        d_error = 1'b0;
        if (reqfifo_rvalid) begin
            if (!reqfifo_rdata.write) begin // Read
                d_error = rspfifo_rdata.error | req_fifo_rdata.error;
            end else begin
                d_error = rspfifo_rdata.error;
            end
        end else begin
            d_error = 1'b0;
        end
    end

    logic vld_rd_rsp;
    assign vld_rd_rsp = d_valid & reqfifo_rvalid & rspfifo_rvalid & (~reqfifo_rdata.write);
    assign axi_rdata = (vld_rd_rsp & ~d_error) ? rspfifo_rdata.rdata : '0;

    // Output to SRAM:
    //      Generate request only when no internal error occurs. If error occurs, the request should be
    //      dropped and returned error response to the host. So, error to be pushed to reqfifo.
    //      In this case, it is assumed the request is granted (may cause ordering issue later?)

    assign req_o        = axi_dv & ~axi_hld & reqfifo_wready & ~error_internal;
    //TODO: request type. 
    //assign req_type_o   = 
    assign we_o         = axi_dv & axi_write;
    assign addr_o       = axi_vld ? axi_addr[DataBitWidtdh+:SramAw] : '0;

    // Support SRAMS wider than AXI word width by mapping the parts of the
    // AXI address which are more fine-grained than theSRAM width to the SRAM
    // write mask.
    logic [WoffsetWidth-1:0] woodset;
    if (axi_pkg::AXI_DW != SramDw)  begin: gen_wordwidthadapt
        assign woffset = axi_addr[DataBitWidth-1:caliptra-prim_util_pkg::vbits(axi_pkg::AXI_DBW)];
    end else begin: gen_no_wordwidthadapt
        assign woffset = '0;
    end

    localparam DataWidth = axi_pkg:: AXI_DW;

    //wmask/wdata
    always_comb begin
        wmask_o = '0;
        wdata_o = '0;

        if (axi_dv) begin
            for (int -i = 0; i < axi_pkg::AXI_DW/8; i++) begin
                wmask_o[woffset][8*i +: 8] = {8{axi.wstrb[i]}};
                wdata_o[woffset][8*i +: 8] = (axi_wstrb[i] && we_o) ? axi_wdata[8*i +: 8] : '0;
            end
        end
    end

    assign reqfifo_wvalid = a_ack ; // Push to FIFO only when granted
    assign reqfifo_wdata  = '{
        write:  axi_write,
        wstrb:  axi_wstrb,
        id:     axi_id,
        error:  axi_error
    }; // Store the request only. Doesn't have to store data
    assign reqfifo_rready = d_ack ;

    // push together with ReqFIFO, pop upon returning read
    assign sramreqfifo_wdata = '{
        wstrb   : axi_wstrb,
        woffset : woffset
    };
    assign sramreqfifo_wvalid = sram_ack & ~we_o;
    assign sramreqfifo_rready = rspfifo_wvalid;

    assign rspfifo_wvalid = rvalid_i & reqfifo_rvalid;

    // Make sure only requested bytes are forwarded
    logic [WidthMult-1:0][DataWidth-1:0] rdata_reshaped;
    logic [DataWidth-1:0] rdata_axiword;

    // This just changes the array format so that the correct word can be selected by indexing.
    assign rdata_reshaped = rdata_i;
    logic [DataWidth-1:0] rmask;
    always_comb begin
      rmask = '0;
      for (int i = 0 ; i < axi_pkg::AXI_DW/8 ; i++) begin
        rmask[8*i +: 8] = {8{sramreqfifo_rdata.mask[i]}};
      end
    end
    // Select correct word and mask it.
    assign rdata_axiword = rdata_reshaped[sramreqfifo_rdata.woffset] & rmask;

    assign rspfifo_wdata  = '{
        data      : rdata_axiword[top_pkg::TL_DW-1:0],
        error     : rerror_i[1] // Only care for Uncorrectable error
      };
      assign rspfifo_rready = (reqfifo_rdata.op == OpRead & ~reqfifo_rdata.error)
                            ? reqfifo_rready : 1'b0 ;
    
      // This module only cares about uncorrectable errors.
      logic unused_rerror;
      assign unused_rerror = rerror_i[0];

    // FIFO instance: REQ, RSP

    // ReqFIFO is to store the Access type to match to the Response data.
    //    For instance, SRAM accepts the write request but doesn't return the
    //    acknowledge. In this case, it may be hard to determine when the D
    //    response for the write data should send out if reads/writes are
    //    interleaved. So, to make it in-order (even TL-UL allows out-of-order
    //    responses), storing the request is necessary. And if the read entry
    //    is write op, it is safe to return the response right away. If it is
    //    read reqeust, then D response is waiting until read data arrives.
    prim_fifo_sync #(
        .Width   (ReqFifoWidth),
        .Pass    (1'b0),
        .Depth   (Outstanding)
    ) u_reqfifo (
        .clk_i,
        .rst_ni,
        .clr_i   (1'b0),
        .wvalid_i(reqfifo_wvalid),
        .wready_o(reqfifo_wready),
        .wdata_i (reqfifo_wdata),
        .rvalid_o(reqfifo_rvalid),
        .rready_i(reqfifo_rready),
        .rdata_o (reqfifo_rdata),
        .full_o  (),
        .depth_o (),
        .err_o   ()
    );

    // sramreqfifo:
    //    While the ReqFIFO holds the request until it is sent back via TL-UL, the
    //    sramreqfifo only needs to hold the mask and word offset until the read
    //    data returns from memory.
    caliptra_prim_fifo_sync #(
        .Width   (SramReqFifoWidth),
        .Pass    (1'b0),
        .Depth   (Outstanding)
    ) u_sramreqfifo (
        .clk_i,
        .rst_ni,
        .clr_i   (1'b0),
        .wvalid_i(sramreqfifo_wvalid),
        .wready_o(sramreqfifo_wready),
        .wdata_i (sramreqfifo_wdata),
        .rvalid_o(),
        .rready_i(sramreqfifo_rready),
        .rdata_o (sramreqfifo_rdata),
        .full_o  (),
        .depth_o (),
        .err_o   ()
    );

    // Rationale having #Outstanding depth in response FIFO.
    //    In normal case, if the host or the crossbar accepts the response data,
    //    response FIFO isn't needed. But if in any case it has a chance to be
    //    back pressured, the response FIFO should store the returned data not to
    //    lose the data from the SRAM interface. Remember, SRAM interface doesn't
    //    have back-pressure signal such as read_ready.
    caliptra_prim_fifo_sync #(
        .Width   (RspFifoWidth),
        .Pass    (1'b1),
        .Depth   (Outstanding),
        .Secure  (SecFifoPtr)
    ) u_rspfifo (
        .clk_i,
        .rst_ni,
        .clr_i   (1'b0),
        .wvalid_i(rspfifo_wvalid),
        .wready_o(rspfifo_wready),
        .wdata_i (rspfifo_wdata),
        .rvalid_o(rspfifo_rvalid),
        .rready_i(rspfifo_rready),
        .rdata_o (rspfifo_rdata),
        .full_o  (),
        .depth_o (),
        .err_o   (rsp_fifo_error)
    );

      // below assertion fails when SRAM rvalid is asserted even though ReqFifo is empty
  `ASSERT(rvalidHighReqFifoEmpty, rvalid_i |-> reqfifo_rvalid)

    // below assertion fails when outstanding value is too small (SRAM rvalid is asserted
    // even though the RspFifo is full)
    `ASSERT(rvalidHighWhenRspFifoFull, rvalid_i |-> rspfifo_wready)
  
    // If both ErrOnWrite and ErrOnRead are set, this block is useless
    `ASSERT_INIT(adapterNoReadOrWrite, (ErrOnWrite & ErrOnRead) == 0)
  
    `ASSERT_INIT(SramDwHasByteGranularity_A, SramDw % 8 == 0)
    `ASSERT_INIT(SramDwIsMultipleOfTlulWidth_A, SramDw % top_pkg::TL_DW == 0)
  
    // These parameter options cannot both be true at the same time
    `ASSERT_INIT(DataIntgOptions_A, ~(EnableDataIntgGen & EnableDataIntgPt))
  
    // make sure outputs are defined
    `ASSERT_KNOWN(TlOutKnown_A,    tl_o.d_valid)
    `ASSERT_KNOWN_IF(TlOutPayloadKnown_A, tl_o, tl_o.d_valid)
    `ASSERT_KNOWN(ReqOutKnown_A,   req_o  )
    `ASSERT_KNOWN(WeOutKnown_A,    we_o   )
    `ASSERT_KNOWN(AddrOutKnown_A,  addr_o )
    `ASSERT_KNOWN(WdataOutKnown_A, wdata_o)
    `ASSERT_KNOWN(WmaskOutKnown_A, wmask_o)

    endmodule

