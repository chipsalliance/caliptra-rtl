../uvm/uvm_reg.sv