// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


module axi_dma_cov_bind;
  `ifdef FCOV
  bind axi_dma_top axi_dma_top_cov_if i_axi_dma_top_cov_if(.*);
  bind axi_dma_top axi_dma_top_cov_props i_axi_dma_top_cov_props(.*);
  `endif
endmodule
