//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.1
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef enum bit[2:0] {reset_op = 3'b000, sha224_op = 3'b100, sha256_op = 3'b101, sha384_op = 3'b110, sha512_op = 3'b111} sha512_in_op_transactions;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

