// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
`ifndef CALIPTRA_REG_DEFINES_HEADER
`define CALIPTRA_REG_DEFINES_HEADER


`define CLP_BASE_ADDR                                                                               (32'h0)
`define CLP_DOE_REG_BASE_ADDR                                                                       (32'h10000000)
`define CLP_DOE_REG_DOE_IV_0                                                                        (32'h10000000)
`define DOE_REG_DOE_IV_0                                                                            (32'h0)
`define CLP_DOE_REG_DOE_IV_1                                                                        (32'h10000004)
`define DOE_REG_DOE_IV_1                                                                            (32'h4)
`define CLP_DOE_REG_DOE_IV_2                                                                        (32'h10000008)
`define DOE_REG_DOE_IV_2                                                                            (32'h8)
`define CLP_DOE_REG_DOE_IV_3                                                                        (32'h1000000c)
`define DOE_REG_DOE_IV_3                                                                            (32'hc)
`define CLP_DOE_REG_DOE_CTRL                                                                        (32'h10000010)
`define DOE_REG_DOE_CTRL                                                                            (32'h10)
`define DOE_REG_DOE_CTRL_CMD_LOW                                                                    (0)
`define DOE_REG_DOE_CTRL_CMD_MASK                                                                   (32'h3)
`define DOE_REG_DOE_CTRL_DEST_LOW                                                                   (2)
`define DOE_REG_DOE_CTRL_DEST_MASK                                                                  (32'h7c)
`define CLP_DOE_REG_DOE_STATUS                                                                      (32'h10000014)
`define DOE_REG_DOE_STATUS                                                                          (32'h14)
`define DOE_REG_DOE_STATUS_READY_LOW                                                                (0)
`define DOE_REG_DOE_STATUS_READY_MASK                                                               (32'h1)
`define DOE_REG_DOE_STATUS_VALID_LOW                                                                (1)
`define DOE_REG_DOE_STATUS_VALID_MASK                                                               (32'h2)
`define DOE_REG_DOE_STATUS_UDS_FLOW_DONE_LOW                                                        (2)
`define DOE_REG_DOE_STATUS_UDS_FLOW_DONE_MASK                                                       (32'h4)
`define DOE_REG_DOE_STATUS_FE_FLOW_DONE_LOW                                                         (3)
`define DOE_REG_DOE_STATUS_FE_FLOW_DONE_MASK                                                        (32'h8)
`define DOE_REG_DOE_STATUS_DEOBF_SECRETS_CLEARED_LOW                                                (4)
`define DOE_REG_DOE_STATUS_DEOBF_SECRETS_CLEARED_MASK                                               (32'h10)
`define CLP_DOE_REG_INTR_BLOCK_RF_START                                                             (32'h10000800)
`define CLP_DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10000800)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                      (32'h800)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                         (0)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                        (32'h1)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                         (1)
`define DOE_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                        (32'h2)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10000804)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                       (32'h804)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                         (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                        (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                         (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                        (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                         (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                        (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                         (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                        (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10000808)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                       (32'h808)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                 (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                                (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1000080c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                   (32'h80c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10000810)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                   (32'h810)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10000814)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                 (32'h814)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                                  (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                                 (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                                  (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                                 (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                                  (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                                 (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                                  (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                                 (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10000818)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                 (32'h818)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                          (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                         (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1000081c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                     (32'h81c)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                     (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                    (32'h1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                     (1)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                    (32'h2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                     (2)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                    (32'h4)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                     (3)
`define DOE_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                    (32'h8)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10000820)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                     (32'h820)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                             (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                            (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                               (32'h10000900)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                   (32'h900)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                               (32'h10000904)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                   (32'h904)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                               (32'h10000908)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                   (32'h908)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                               (32'h1000090c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                   (32'h90c)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10000980)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                           (32'h980)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                          (32'h10000a00)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                              (32'ha00)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                          (32'h10000a04)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                              (32'ha04)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                          (32'h10000a08)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                              (32'ha08)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                          (32'h10000a0c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                              (32'ha0c)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                    (0)
`define DOE_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                   (32'h1)
`define CLP_DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10000a10)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                      (32'ha10)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define DOE_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_ECC_REG_BASE_ADDR                                                                       (32'h10008000)
`define CLP_ECC_REG_ECC_NAME_0                                                                      (32'h10008000)
`define ECC_REG_ECC_NAME_0                                                                          (32'h0)
`define CLP_ECC_REG_ECC_NAME_1                                                                      (32'h10008004)
`define ECC_REG_ECC_NAME_1                                                                          (32'h4)
`define CLP_ECC_REG_ECC_VERSION_0                                                                   (32'h10008008)
`define ECC_REG_ECC_VERSION_0                                                                       (32'h8)
`define CLP_ECC_REG_ECC_VERSION_1                                                                   (32'h1000800c)
`define ECC_REG_ECC_VERSION_1                                                                       (32'hc)
`define CLP_ECC_REG_ECC_CTRL                                                                        (32'h10008010)
`define ECC_REG_ECC_CTRL                                                                            (32'h10)
`define ECC_REG_ECC_CTRL_CTRL_LOW                                                                   (0)
`define ECC_REG_ECC_CTRL_CTRL_MASK                                                                  (32'h3)
`define ECC_REG_ECC_CTRL_ZEROIZE_LOW                                                                (2)
`define ECC_REG_ECC_CTRL_ZEROIZE_MASK                                                               (32'h4)
`define ECC_REG_ECC_CTRL_PCR_SIGN_LOW                                                               (3)
`define ECC_REG_ECC_CTRL_PCR_SIGN_MASK                                                              (32'h8)
`define CLP_ECC_REG_ECC_STATUS                                                                      (32'h10008018)
`define ECC_REG_ECC_STATUS                                                                          (32'h18)
`define ECC_REG_ECC_STATUS_READY_LOW                                                                (0)
`define ECC_REG_ECC_STATUS_READY_MASK                                                               (32'h1)
`define ECC_REG_ECC_STATUS_VALID_LOW                                                                (1)
`define ECC_REG_ECC_STATUS_VALID_MASK                                                               (32'h2)
`define CLP_ECC_REG_ECC_SCACONFIG                                                                   (32'h10008020)
`define ECC_REG_ECC_SCACONFIG                                                                       (32'h20)
`define ECC_REG_ECC_SCACONFIG_POINT_RND_EN_LOW                                                      (0)
`define ECC_REG_ECC_SCACONFIG_POINT_RND_EN_MASK                                                     (32'h1)
`define ECC_REG_ECC_SCACONFIG_MASK_SIGN_EN_LOW                                                      (1)
`define ECC_REG_ECC_SCACONFIG_MASK_SIGN_EN_MASK                                                     (32'h2)
`define ECC_REG_ECC_SCACONFIG_SCALAR_RND_EN_LOW                                                     (2)
`define ECC_REG_ECC_SCACONFIG_SCALAR_RND_EN_MASK                                                    (32'h4)
`define CLP_ECC_REG_ECC_SEED_0                                                                      (32'h10008080)
`define ECC_REG_ECC_SEED_0                                                                          (32'h80)
`define CLP_ECC_REG_ECC_SEED_1                                                                      (32'h10008084)
`define ECC_REG_ECC_SEED_1                                                                          (32'h84)
`define CLP_ECC_REG_ECC_SEED_2                                                                      (32'h10008088)
`define ECC_REG_ECC_SEED_2                                                                          (32'h88)
`define CLP_ECC_REG_ECC_SEED_3                                                                      (32'h1000808c)
`define ECC_REG_ECC_SEED_3                                                                          (32'h8c)
`define CLP_ECC_REG_ECC_SEED_4                                                                      (32'h10008090)
`define ECC_REG_ECC_SEED_4                                                                          (32'h90)
`define CLP_ECC_REG_ECC_SEED_5                                                                      (32'h10008094)
`define ECC_REG_ECC_SEED_5                                                                          (32'h94)
`define CLP_ECC_REG_ECC_SEED_6                                                                      (32'h10008098)
`define ECC_REG_ECC_SEED_6                                                                          (32'h98)
`define CLP_ECC_REG_ECC_SEED_7                                                                      (32'h1000809c)
`define ECC_REG_ECC_SEED_7                                                                          (32'h9c)
`define CLP_ECC_REG_ECC_SEED_8                                                                      (32'h100080a0)
`define ECC_REG_ECC_SEED_8                                                                          (32'ha0)
`define CLP_ECC_REG_ECC_SEED_9                                                                      (32'h100080a4)
`define ECC_REG_ECC_SEED_9                                                                          (32'ha4)
`define CLP_ECC_REG_ECC_SEED_10                                                                     (32'h100080a8)
`define ECC_REG_ECC_SEED_10                                                                         (32'ha8)
`define CLP_ECC_REG_ECC_SEED_11                                                                     (32'h100080ac)
`define ECC_REG_ECC_SEED_11                                                                         (32'hac)
`define CLP_ECC_REG_ECC_MSG_0                                                                       (32'h10008100)
`define ECC_REG_ECC_MSG_0                                                                           (32'h100)
`define CLP_ECC_REG_ECC_MSG_1                                                                       (32'h10008104)
`define ECC_REG_ECC_MSG_1                                                                           (32'h104)
`define CLP_ECC_REG_ECC_MSG_2                                                                       (32'h10008108)
`define ECC_REG_ECC_MSG_2                                                                           (32'h108)
`define CLP_ECC_REG_ECC_MSG_3                                                                       (32'h1000810c)
`define ECC_REG_ECC_MSG_3                                                                           (32'h10c)
`define CLP_ECC_REG_ECC_MSG_4                                                                       (32'h10008110)
`define ECC_REG_ECC_MSG_4                                                                           (32'h110)
`define CLP_ECC_REG_ECC_MSG_5                                                                       (32'h10008114)
`define ECC_REG_ECC_MSG_5                                                                           (32'h114)
`define CLP_ECC_REG_ECC_MSG_6                                                                       (32'h10008118)
`define ECC_REG_ECC_MSG_6                                                                           (32'h118)
`define CLP_ECC_REG_ECC_MSG_7                                                                       (32'h1000811c)
`define ECC_REG_ECC_MSG_7                                                                           (32'h11c)
`define CLP_ECC_REG_ECC_MSG_8                                                                       (32'h10008120)
`define ECC_REG_ECC_MSG_8                                                                           (32'h120)
`define CLP_ECC_REG_ECC_MSG_9                                                                       (32'h10008124)
`define ECC_REG_ECC_MSG_9                                                                           (32'h124)
`define CLP_ECC_REG_ECC_MSG_10                                                                      (32'h10008128)
`define ECC_REG_ECC_MSG_10                                                                          (32'h128)
`define CLP_ECC_REG_ECC_MSG_11                                                                      (32'h1000812c)
`define ECC_REG_ECC_MSG_11                                                                          (32'h12c)
`define CLP_ECC_REG_ECC_PRIVKEY_0                                                                   (32'h10008180)
`define ECC_REG_ECC_PRIVKEY_0                                                                       (32'h180)
`define CLP_ECC_REG_ECC_PRIVKEY_1                                                                   (32'h10008184)
`define ECC_REG_ECC_PRIVKEY_1                                                                       (32'h184)
`define CLP_ECC_REG_ECC_PRIVKEY_2                                                                   (32'h10008188)
`define ECC_REG_ECC_PRIVKEY_2                                                                       (32'h188)
`define CLP_ECC_REG_ECC_PRIVKEY_3                                                                   (32'h1000818c)
`define ECC_REG_ECC_PRIVKEY_3                                                                       (32'h18c)
`define CLP_ECC_REG_ECC_PRIVKEY_4                                                                   (32'h10008190)
`define ECC_REG_ECC_PRIVKEY_4                                                                       (32'h190)
`define CLP_ECC_REG_ECC_PRIVKEY_5                                                                   (32'h10008194)
`define ECC_REG_ECC_PRIVKEY_5                                                                       (32'h194)
`define CLP_ECC_REG_ECC_PRIVKEY_6                                                                   (32'h10008198)
`define ECC_REG_ECC_PRIVKEY_6                                                                       (32'h198)
`define CLP_ECC_REG_ECC_PRIVKEY_7                                                                   (32'h1000819c)
`define ECC_REG_ECC_PRIVKEY_7                                                                       (32'h19c)
`define CLP_ECC_REG_ECC_PRIVKEY_8                                                                   (32'h100081a0)
`define ECC_REG_ECC_PRIVKEY_8                                                                       (32'h1a0)
`define CLP_ECC_REG_ECC_PRIVKEY_9                                                                   (32'h100081a4)
`define ECC_REG_ECC_PRIVKEY_9                                                                       (32'h1a4)
`define CLP_ECC_REG_ECC_PRIVKEY_10                                                                  (32'h100081a8)
`define ECC_REG_ECC_PRIVKEY_10                                                                      (32'h1a8)
`define CLP_ECC_REG_ECC_PRIVKEY_11                                                                  (32'h100081ac)
`define ECC_REG_ECC_PRIVKEY_11                                                                      (32'h1ac)
`define CLP_ECC_REG_ECC_PUBKEY_X_0                                                                  (32'h10008200)
`define ECC_REG_ECC_PUBKEY_X_0                                                                      (32'h200)
`define CLP_ECC_REG_ECC_PUBKEY_X_1                                                                  (32'h10008204)
`define ECC_REG_ECC_PUBKEY_X_1                                                                      (32'h204)
`define CLP_ECC_REG_ECC_PUBKEY_X_2                                                                  (32'h10008208)
`define ECC_REG_ECC_PUBKEY_X_2                                                                      (32'h208)
`define CLP_ECC_REG_ECC_PUBKEY_X_3                                                                  (32'h1000820c)
`define ECC_REG_ECC_PUBKEY_X_3                                                                      (32'h20c)
`define CLP_ECC_REG_ECC_PUBKEY_X_4                                                                  (32'h10008210)
`define ECC_REG_ECC_PUBKEY_X_4                                                                      (32'h210)
`define CLP_ECC_REG_ECC_PUBKEY_X_5                                                                  (32'h10008214)
`define ECC_REG_ECC_PUBKEY_X_5                                                                      (32'h214)
`define CLP_ECC_REG_ECC_PUBKEY_X_6                                                                  (32'h10008218)
`define ECC_REG_ECC_PUBKEY_X_6                                                                      (32'h218)
`define CLP_ECC_REG_ECC_PUBKEY_X_7                                                                  (32'h1000821c)
`define ECC_REG_ECC_PUBKEY_X_7                                                                      (32'h21c)
`define CLP_ECC_REG_ECC_PUBKEY_X_8                                                                  (32'h10008220)
`define ECC_REG_ECC_PUBKEY_X_8                                                                      (32'h220)
`define CLP_ECC_REG_ECC_PUBKEY_X_9                                                                  (32'h10008224)
`define ECC_REG_ECC_PUBKEY_X_9                                                                      (32'h224)
`define CLP_ECC_REG_ECC_PUBKEY_X_10                                                                 (32'h10008228)
`define ECC_REG_ECC_PUBKEY_X_10                                                                     (32'h228)
`define CLP_ECC_REG_ECC_PUBKEY_X_11                                                                 (32'h1000822c)
`define ECC_REG_ECC_PUBKEY_X_11                                                                     (32'h22c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_0                                                                  (32'h10008280)
`define ECC_REG_ECC_PUBKEY_Y_0                                                                      (32'h280)
`define CLP_ECC_REG_ECC_PUBKEY_Y_1                                                                  (32'h10008284)
`define ECC_REG_ECC_PUBKEY_Y_1                                                                      (32'h284)
`define CLP_ECC_REG_ECC_PUBKEY_Y_2                                                                  (32'h10008288)
`define ECC_REG_ECC_PUBKEY_Y_2                                                                      (32'h288)
`define CLP_ECC_REG_ECC_PUBKEY_Y_3                                                                  (32'h1000828c)
`define ECC_REG_ECC_PUBKEY_Y_3                                                                      (32'h28c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_4                                                                  (32'h10008290)
`define ECC_REG_ECC_PUBKEY_Y_4                                                                      (32'h290)
`define CLP_ECC_REG_ECC_PUBKEY_Y_5                                                                  (32'h10008294)
`define ECC_REG_ECC_PUBKEY_Y_5                                                                      (32'h294)
`define CLP_ECC_REG_ECC_PUBKEY_Y_6                                                                  (32'h10008298)
`define ECC_REG_ECC_PUBKEY_Y_6                                                                      (32'h298)
`define CLP_ECC_REG_ECC_PUBKEY_Y_7                                                                  (32'h1000829c)
`define ECC_REG_ECC_PUBKEY_Y_7                                                                      (32'h29c)
`define CLP_ECC_REG_ECC_PUBKEY_Y_8                                                                  (32'h100082a0)
`define ECC_REG_ECC_PUBKEY_Y_8                                                                      (32'h2a0)
`define CLP_ECC_REG_ECC_PUBKEY_Y_9                                                                  (32'h100082a4)
`define ECC_REG_ECC_PUBKEY_Y_9                                                                      (32'h2a4)
`define CLP_ECC_REG_ECC_PUBKEY_Y_10                                                                 (32'h100082a8)
`define ECC_REG_ECC_PUBKEY_Y_10                                                                     (32'h2a8)
`define CLP_ECC_REG_ECC_PUBKEY_Y_11                                                                 (32'h100082ac)
`define ECC_REG_ECC_PUBKEY_Y_11                                                                     (32'h2ac)
`define CLP_ECC_REG_ECC_SIGN_R_0                                                                    (32'h10008300)
`define ECC_REG_ECC_SIGN_R_0                                                                        (32'h300)
`define CLP_ECC_REG_ECC_SIGN_R_1                                                                    (32'h10008304)
`define ECC_REG_ECC_SIGN_R_1                                                                        (32'h304)
`define CLP_ECC_REG_ECC_SIGN_R_2                                                                    (32'h10008308)
`define ECC_REG_ECC_SIGN_R_2                                                                        (32'h308)
`define CLP_ECC_REG_ECC_SIGN_R_3                                                                    (32'h1000830c)
`define ECC_REG_ECC_SIGN_R_3                                                                        (32'h30c)
`define CLP_ECC_REG_ECC_SIGN_R_4                                                                    (32'h10008310)
`define ECC_REG_ECC_SIGN_R_4                                                                        (32'h310)
`define CLP_ECC_REG_ECC_SIGN_R_5                                                                    (32'h10008314)
`define ECC_REG_ECC_SIGN_R_5                                                                        (32'h314)
`define CLP_ECC_REG_ECC_SIGN_R_6                                                                    (32'h10008318)
`define ECC_REG_ECC_SIGN_R_6                                                                        (32'h318)
`define CLP_ECC_REG_ECC_SIGN_R_7                                                                    (32'h1000831c)
`define ECC_REG_ECC_SIGN_R_7                                                                        (32'h31c)
`define CLP_ECC_REG_ECC_SIGN_R_8                                                                    (32'h10008320)
`define ECC_REG_ECC_SIGN_R_8                                                                        (32'h320)
`define CLP_ECC_REG_ECC_SIGN_R_9                                                                    (32'h10008324)
`define ECC_REG_ECC_SIGN_R_9                                                                        (32'h324)
`define CLP_ECC_REG_ECC_SIGN_R_10                                                                   (32'h10008328)
`define ECC_REG_ECC_SIGN_R_10                                                                       (32'h328)
`define CLP_ECC_REG_ECC_SIGN_R_11                                                                   (32'h1000832c)
`define ECC_REG_ECC_SIGN_R_11                                                                       (32'h32c)
`define CLP_ECC_REG_ECC_SIGN_S_0                                                                    (32'h10008380)
`define ECC_REG_ECC_SIGN_S_0                                                                        (32'h380)
`define CLP_ECC_REG_ECC_SIGN_S_1                                                                    (32'h10008384)
`define ECC_REG_ECC_SIGN_S_1                                                                        (32'h384)
`define CLP_ECC_REG_ECC_SIGN_S_2                                                                    (32'h10008388)
`define ECC_REG_ECC_SIGN_S_2                                                                        (32'h388)
`define CLP_ECC_REG_ECC_SIGN_S_3                                                                    (32'h1000838c)
`define ECC_REG_ECC_SIGN_S_3                                                                        (32'h38c)
`define CLP_ECC_REG_ECC_SIGN_S_4                                                                    (32'h10008390)
`define ECC_REG_ECC_SIGN_S_4                                                                        (32'h390)
`define CLP_ECC_REG_ECC_SIGN_S_5                                                                    (32'h10008394)
`define ECC_REG_ECC_SIGN_S_5                                                                        (32'h394)
`define CLP_ECC_REG_ECC_SIGN_S_6                                                                    (32'h10008398)
`define ECC_REG_ECC_SIGN_S_6                                                                        (32'h398)
`define CLP_ECC_REG_ECC_SIGN_S_7                                                                    (32'h1000839c)
`define ECC_REG_ECC_SIGN_S_7                                                                        (32'h39c)
`define CLP_ECC_REG_ECC_SIGN_S_8                                                                    (32'h100083a0)
`define ECC_REG_ECC_SIGN_S_8                                                                        (32'h3a0)
`define CLP_ECC_REG_ECC_SIGN_S_9                                                                    (32'h100083a4)
`define ECC_REG_ECC_SIGN_S_9                                                                        (32'h3a4)
`define CLP_ECC_REG_ECC_SIGN_S_10                                                                   (32'h100083a8)
`define ECC_REG_ECC_SIGN_S_10                                                                       (32'h3a8)
`define CLP_ECC_REG_ECC_SIGN_S_11                                                                   (32'h100083ac)
`define ECC_REG_ECC_SIGN_S_11                                                                       (32'h3ac)
`define CLP_ECC_REG_ECC_VERIFY_R_0                                                                  (32'h10008400)
`define ECC_REG_ECC_VERIFY_R_0                                                                      (32'h400)
`define CLP_ECC_REG_ECC_VERIFY_R_1                                                                  (32'h10008404)
`define ECC_REG_ECC_VERIFY_R_1                                                                      (32'h404)
`define CLP_ECC_REG_ECC_VERIFY_R_2                                                                  (32'h10008408)
`define ECC_REG_ECC_VERIFY_R_2                                                                      (32'h408)
`define CLP_ECC_REG_ECC_VERIFY_R_3                                                                  (32'h1000840c)
`define ECC_REG_ECC_VERIFY_R_3                                                                      (32'h40c)
`define CLP_ECC_REG_ECC_VERIFY_R_4                                                                  (32'h10008410)
`define ECC_REG_ECC_VERIFY_R_4                                                                      (32'h410)
`define CLP_ECC_REG_ECC_VERIFY_R_5                                                                  (32'h10008414)
`define ECC_REG_ECC_VERIFY_R_5                                                                      (32'h414)
`define CLP_ECC_REG_ECC_VERIFY_R_6                                                                  (32'h10008418)
`define ECC_REG_ECC_VERIFY_R_6                                                                      (32'h418)
`define CLP_ECC_REG_ECC_VERIFY_R_7                                                                  (32'h1000841c)
`define ECC_REG_ECC_VERIFY_R_7                                                                      (32'h41c)
`define CLP_ECC_REG_ECC_VERIFY_R_8                                                                  (32'h10008420)
`define ECC_REG_ECC_VERIFY_R_8                                                                      (32'h420)
`define CLP_ECC_REG_ECC_VERIFY_R_9                                                                  (32'h10008424)
`define ECC_REG_ECC_VERIFY_R_9                                                                      (32'h424)
`define CLP_ECC_REG_ECC_VERIFY_R_10                                                                 (32'h10008428)
`define ECC_REG_ECC_VERIFY_R_10                                                                     (32'h428)
`define CLP_ECC_REG_ECC_VERIFY_R_11                                                                 (32'h1000842c)
`define ECC_REG_ECC_VERIFY_R_11                                                                     (32'h42c)
`define CLP_ECC_REG_ECC_IV_0                                                                        (32'h10008480)
`define ECC_REG_ECC_IV_0                                                                            (32'h480)
`define CLP_ECC_REG_ECC_IV_1                                                                        (32'h10008484)
`define ECC_REG_ECC_IV_1                                                                            (32'h484)
`define CLP_ECC_REG_ECC_IV_2                                                                        (32'h10008488)
`define ECC_REG_ECC_IV_2                                                                            (32'h488)
`define CLP_ECC_REG_ECC_IV_3                                                                        (32'h1000848c)
`define ECC_REG_ECC_IV_3                                                                            (32'h48c)
`define CLP_ECC_REG_ECC_IV_4                                                                        (32'h10008490)
`define ECC_REG_ECC_IV_4                                                                            (32'h490)
`define CLP_ECC_REG_ECC_IV_5                                                                        (32'h10008494)
`define ECC_REG_ECC_IV_5                                                                            (32'h494)
`define CLP_ECC_REG_ECC_IV_6                                                                        (32'h10008498)
`define ECC_REG_ECC_IV_6                                                                            (32'h498)
`define CLP_ECC_REG_ECC_IV_7                                                                        (32'h1000849c)
`define ECC_REG_ECC_IV_7                                                                            (32'h49c)
`define CLP_ECC_REG_ECC_IV_8                                                                        (32'h100084a0)
`define ECC_REG_ECC_IV_8                                                                            (32'h4a0)
`define CLP_ECC_REG_ECC_IV_9                                                                        (32'h100084a4)
`define ECC_REG_ECC_IV_9                                                                            (32'h4a4)
`define CLP_ECC_REG_ECC_IV_10                                                                       (32'h100084a8)
`define ECC_REG_ECC_IV_10                                                                           (32'h4a8)
`define CLP_ECC_REG_ECC_IV_11                                                                       (32'h100084ac)
`define ECC_REG_ECC_IV_11                                                                           (32'h4ac)
`define CLP_ECC_REG_ECC_NONCE_0                                                                     (32'h10008500)
`define ECC_REG_ECC_NONCE_0                                                                         (32'h500)
`define CLP_ECC_REG_ECC_NONCE_1                                                                     (32'h10008504)
`define ECC_REG_ECC_NONCE_1                                                                         (32'h504)
`define CLP_ECC_REG_ECC_NONCE_2                                                                     (32'h10008508)
`define ECC_REG_ECC_NONCE_2                                                                         (32'h508)
`define CLP_ECC_REG_ECC_NONCE_3                                                                     (32'h1000850c)
`define ECC_REG_ECC_NONCE_3                                                                         (32'h50c)
`define CLP_ECC_REG_ECC_NONCE_4                                                                     (32'h10008510)
`define ECC_REG_ECC_NONCE_4                                                                         (32'h510)
`define CLP_ECC_REG_ECC_NONCE_5                                                                     (32'h10008514)
`define ECC_REG_ECC_NONCE_5                                                                         (32'h514)
`define CLP_ECC_REG_ECC_NONCE_6                                                                     (32'h10008518)
`define ECC_REG_ECC_NONCE_6                                                                         (32'h518)
`define CLP_ECC_REG_ECC_NONCE_7                                                                     (32'h1000851c)
`define ECC_REG_ECC_NONCE_7                                                                         (32'h51c)
`define CLP_ECC_REG_ECC_NONCE_8                                                                     (32'h10008520)
`define ECC_REG_ECC_NONCE_8                                                                         (32'h520)
`define CLP_ECC_REG_ECC_NONCE_9                                                                     (32'h10008524)
`define ECC_REG_ECC_NONCE_9                                                                         (32'h524)
`define CLP_ECC_REG_ECC_NONCE_10                                                                    (32'h10008528)
`define ECC_REG_ECC_NONCE_10                                                                        (32'h528)
`define CLP_ECC_REG_ECC_NONCE_11                                                                    (32'h1000852c)
`define ECC_REG_ECC_NONCE_11                                                                        (32'h52c)
`define CLP_ECC_REG_ECC_KV_RD_PKEY_CTRL                                                             (32'h10008600)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL                                                                 (32'h600)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_EN_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_EN_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_ENTRY_LOW                                                  (1)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_READ_ENTRY_MASK                                                 (32'h3e)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_PCR_HASH_EXTEND_LOW                                             (6)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_PCR_HASH_EXTEND_MASK                                            (32'h40)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_RSVD_LOW                                                        (7)
`define ECC_REG_ECC_KV_RD_PKEY_CTRL_RSVD_MASK                                                       (32'hffffff80)
`define CLP_ECC_REG_ECC_KV_RD_PKEY_STATUS                                                           (32'h10008604)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS                                                               (32'h604)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_RD_PKEY_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_ECC_KV_RD_SEED_CTRL                                                             (32'h10008608)
`define ECC_REG_ECC_KV_RD_SEED_CTRL                                                                 (32'h608)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_EN_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_EN_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_ENTRY_LOW                                                  (1)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_READ_ENTRY_MASK                                                 (32'h3e)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_PCR_HASH_EXTEND_LOW                                             (6)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_PCR_HASH_EXTEND_MASK                                            (32'h40)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_RSVD_LOW                                                        (7)
`define ECC_REG_ECC_KV_RD_SEED_CTRL_RSVD_MASK                                                       (32'hffffff80)
`define CLP_ECC_REG_ECC_KV_RD_SEED_STATUS                                                           (32'h1000860c)
`define ECC_REG_ECC_KV_RD_SEED_STATUS                                                               (32'h60c)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_RD_SEED_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_ECC_KV_RD_MSG_CTRL                                                              (32'h10008610)
`define ECC_REG_ECC_KV_RD_MSG_CTRL                                                                  (32'h610)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_READ_EN_LOW                                                      (0)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_READ_EN_MASK                                                     (32'h1)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_READ_ENTRY_LOW                                                   (1)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_READ_ENTRY_MASK                                                  (32'h3e)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_PCR_HASH_EXTEND_LOW                                              (6)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_PCR_HASH_EXTEND_MASK                                             (32'h40)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_RSVD_LOW                                                         (7)
`define ECC_REG_ECC_KV_RD_MSG_CTRL_RSVD_MASK                                                        (32'hffffff80)
`define CLP_ECC_REG_ECC_KV_RD_MSG_STATUS                                                            (32'h10008614)
`define ECC_REG_ECC_KV_RD_MSG_STATUS                                                                (32'h614)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_READY_LOW                                                      (0)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_READY_MASK                                                     (32'h1)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_VALID_LOW                                                      (1)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_VALID_MASK                                                     (32'h2)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_ERROR_LOW                                                      (2)
`define ECC_REG_ECC_KV_RD_MSG_STATUS_ERROR_MASK                                                     (32'h3fc)
`define CLP_ECC_REG_ECC_KV_WR_PKEY_CTRL                                                             (32'h10008618)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL                                                                 (32'h618)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_EN_LOW                                                    (0)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_EN_MASK                                                   (32'h1)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_ENTRY_LOW                                                 (1)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_WRITE_ENTRY_MASK                                                (32'h3e)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_KEY_DEST_VALID_LOW                                         (6)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_KEY_DEST_VALID_MASK                                        (32'h40)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                       (7)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                      (32'h80)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_SHA_BLOCK_DEST_VALID_LOW                                        (8)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_SHA_BLOCK_DEST_VALID_MASK                                       (32'h100)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_PKEY_DEST_VALID_LOW                                         (9)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_PKEY_DEST_VALID_MASK                                        (32'h200)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_SEED_DEST_VALID_LOW                                         (10)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_SEED_DEST_VALID_MASK                                        (32'h400)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_MSG_DEST_VALID_LOW                                          (11)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_ECC_MSG_DEST_VALID_MASK                                         (32'h800)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_RSVD_LOW                                                        (12)
`define ECC_REG_ECC_KV_WR_PKEY_CTRL_RSVD_MASK                                                       (32'hfffff000)
`define CLP_ECC_REG_ECC_KV_WR_PKEY_STATUS                                                           (32'h1000861c)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS                                                               (32'h61c)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_READY_LOW                                                     (0)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_READY_MASK                                                    (32'h1)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_VALID_LOW                                                     (1)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_VALID_MASK                                                    (32'h2)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_ERROR_LOW                                                     (2)
`define ECC_REG_ECC_KV_WR_PKEY_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_ECC_REG_INTR_BLOCK_RF_START                                                             (32'h10008800)
`define CLP_ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h10008800)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                      (32'h800)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                         (0)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                        (32'h1)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                         (1)
`define ECC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                        (32'h2)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h10008804)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                       (32'h804)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_LOW                                 (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_MASK                                (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h10008808)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                       (32'h808)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                 (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                                (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h1000880c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                   (32'h80c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h10008810)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                   (32'h810)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                       (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                      (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h10008814)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                 (32'h814)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_LOW                          (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_MASK                         (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h10008818)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                 (32'h818)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                          (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                         (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h1000881c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                     (32'h81c)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_LOW                             (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_MASK                            (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h10008820)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                     (32'h820)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                             (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                            (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h10008900)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                           (32'h900)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                       (32'h10008980)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                           (32'h980)
`define CLP_ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'h10008a00)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                      (32'ha00)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define ECC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                  (32'h10008a04)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                      (32'ha04)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                            (0)
`define ECC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                           (32'h1)
`define CLP_HMAC_REG_BASE_ADDR                                                                      (32'h10010000)
`define CLP_HMAC_REG_HMAC384_NAME_0                                                                 (32'h10010000)
`define HMAC_REG_HMAC384_NAME_0                                                                     (32'h0)
`define CLP_HMAC_REG_HMAC384_NAME_1                                                                 (32'h10010004)
`define HMAC_REG_HMAC384_NAME_1                                                                     (32'h4)
`define CLP_HMAC_REG_HMAC384_VERSION_0                                                              (32'h10010008)
`define HMAC_REG_HMAC384_VERSION_0                                                                  (32'h8)
`define CLP_HMAC_REG_HMAC384_VERSION_1                                                              (32'h1001000c)
`define HMAC_REG_HMAC384_VERSION_1                                                                  (32'hc)
`define CLP_HMAC_REG_HMAC384_CTRL                                                                   (32'h10010010)
`define HMAC_REG_HMAC384_CTRL                                                                       (32'h10)
`define HMAC_REG_HMAC384_CTRL_INIT_LOW                                                              (0)
`define HMAC_REG_HMAC384_CTRL_INIT_MASK                                                             (32'h1)
`define HMAC_REG_HMAC384_CTRL_NEXT_LOW                                                              (1)
`define HMAC_REG_HMAC384_CTRL_NEXT_MASK                                                             (32'h2)
`define HMAC_REG_HMAC384_CTRL_ZEROIZE_LOW                                                           (2)
`define HMAC_REG_HMAC384_CTRL_ZEROIZE_MASK                                                          (32'h4)
`define CLP_HMAC_REG_HMAC384_STATUS                                                                 (32'h10010018)
`define HMAC_REG_HMAC384_STATUS                                                                     (32'h18)
`define HMAC_REG_HMAC384_STATUS_READY_LOW                                                           (0)
`define HMAC_REG_HMAC384_STATUS_READY_MASK                                                          (32'h1)
`define HMAC_REG_HMAC384_STATUS_VALID_LOW                                                           (1)
`define HMAC_REG_HMAC384_STATUS_VALID_MASK                                                          (32'h2)
`define CLP_HMAC_REG_HMAC384_KEY_0                                                                  (32'h10010040)
`define HMAC_REG_HMAC384_KEY_0                                                                      (32'h40)
`define CLP_HMAC_REG_HMAC384_KEY_1                                                                  (32'h10010044)
`define HMAC_REG_HMAC384_KEY_1                                                                      (32'h44)
`define CLP_HMAC_REG_HMAC384_KEY_2                                                                  (32'h10010048)
`define HMAC_REG_HMAC384_KEY_2                                                                      (32'h48)
`define CLP_HMAC_REG_HMAC384_KEY_3                                                                  (32'h1001004c)
`define HMAC_REG_HMAC384_KEY_3                                                                      (32'h4c)
`define CLP_HMAC_REG_HMAC384_KEY_4                                                                  (32'h10010050)
`define HMAC_REG_HMAC384_KEY_4                                                                      (32'h50)
`define CLP_HMAC_REG_HMAC384_KEY_5                                                                  (32'h10010054)
`define HMAC_REG_HMAC384_KEY_5                                                                      (32'h54)
`define CLP_HMAC_REG_HMAC384_KEY_6                                                                  (32'h10010058)
`define HMAC_REG_HMAC384_KEY_6                                                                      (32'h58)
`define CLP_HMAC_REG_HMAC384_KEY_7                                                                  (32'h1001005c)
`define HMAC_REG_HMAC384_KEY_7                                                                      (32'h5c)
`define CLP_HMAC_REG_HMAC384_KEY_8                                                                  (32'h10010060)
`define HMAC_REG_HMAC384_KEY_8                                                                      (32'h60)
`define CLP_HMAC_REG_HMAC384_KEY_9                                                                  (32'h10010064)
`define HMAC_REG_HMAC384_KEY_9                                                                      (32'h64)
`define CLP_HMAC_REG_HMAC384_KEY_10                                                                 (32'h10010068)
`define HMAC_REG_HMAC384_KEY_10                                                                     (32'h68)
`define CLP_HMAC_REG_HMAC384_KEY_11                                                                 (32'h1001006c)
`define HMAC_REG_HMAC384_KEY_11                                                                     (32'h6c)
`define CLP_HMAC_REG_HMAC384_BLOCK_0                                                                (32'h10010080)
`define HMAC_REG_HMAC384_BLOCK_0                                                                    (32'h80)
`define CLP_HMAC_REG_HMAC384_BLOCK_1                                                                (32'h10010084)
`define HMAC_REG_HMAC384_BLOCK_1                                                                    (32'h84)
`define CLP_HMAC_REG_HMAC384_BLOCK_2                                                                (32'h10010088)
`define HMAC_REG_HMAC384_BLOCK_2                                                                    (32'h88)
`define CLP_HMAC_REG_HMAC384_BLOCK_3                                                                (32'h1001008c)
`define HMAC_REG_HMAC384_BLOCK_3                                                                    (32'h8c)
`define CLP_HMAC_REG_HMAC384_BLOCK_4                                                                (32'h10010090)
`define HMAC_REG_HMAC384_BLOCK_4                                                                    (32'h90)
`define CLP_HMAC_REG_HMAC384_BLOCK_5                                                                (32'h10010094)
`define HMAC_REG_HMAC384_BLOCK_5                                                                    (32'h94)
`define CLP_HMAC_REG_HMAC384_BLOCK_6                                                                (32'h10010098)
`define HMAC_REG_HMAC384_BLOCK_6                                                                    (32'h98)
`define CLP_HMAC_REG_HMAC384_BLOCK_7                                                                (32'h1001009c)
`define HMAC_REG_HMAC384_BLOCK_7                                                                    (32'h9c)
`define CLP_HMAC_REG_HMAC384_BLOCK_8                                                                (32'h100100a0)
`define HMAC_REG_HMAC384_BLOCK_8                                                                    (32'ha0)
`define CLP_HMAC_REG_HMAC384_BLOCK_9                                                                (32'h100100a4)
`define HMAC_REG_HMAC384_BLOCK_9                                                                    (32'ha4)
`define CLP_HMAC_REG_HMAC384_BLOCK_10                                                               (32'h100100a8)
`define HMAC_REG_HMAC384_BLOCK_10                                                                   (32'ha8)
`define CLP_HMAC_REG_HMAC384_BLOCK_11                                                               (32'h100100ac)
`define HMAC_REG_HMAC384_BLOCK_11                                                                   (32'hac)
`define CLP_HMAC_REG_HMAC384_BLOCK_12                                                               (32'h100100b0)
`define HMAC_REG_HMAC384_BLOCK_12                                                                   (32'hb0)
`define CLP_HMAC_REG_HMAC384_BLOCK_13                                                               (32'h100100b4)
`define HMAC_REG_HMAC384_BLOCK_13                                                                   (32'hb4)
`define CLP_HMAC_REG_HMAC384_BLOCK_14                                                               (32'h100100b8)
`define HMAC_REG_HMAC384_BLOCK_14                                                                   (32'hb8)
`define CLP_HMAC_REG_HMAC384_BLOCK_15                                                               (32'h100100bc)
`define HMAC_REG_HMAC384_BLOCK_15                                                                   (32'hbc)
`define CLP_HMAC_REG_HMAC384_BLOCK_16                                                               (32'h100100c0)
`define HMAC_REG_HMAC384_BLOCK_16                                                                   (32'hc0)
`define CLP_HMAC_REG_HMAC384_BLOCK_17                                                               (32'h100100c4)
`define HMAC_REG_HMAC384_BLOCK_17                                                                   (32'hc4)
`define CLP_HMAC_REG_HMAC384_BLOCK_18                                                               (32'h100100c8)
`define HMAC_REG_HMAC384_BLOCK_18                                                                   (32'hc8)
`define CLP_HMAC_REG_HMAC384_BLOCK_19                                                               (32'h100100cc)
`define HMAC_REG_HMAC384_BLOCK_19                                                                   (32'hcc)
`define CLP_HMAC_REG_HMAC384_BLOCK_20                                                               (32'h100100d0)
`define HMAC_REG_HMAC384_BLOCK_20                                                                   (32'hd0)
`define CLP_HMAC_REG_HMAC384_BLOCK_21                                                               (32'h100100d4)
`define HMAC_REG_HMAC384_BLOCK_21                                                                   (32'hd4)
`define CLP_HMAC_REG_HMAC384_BLOCK_22                                                               (32'h100100d8)
`define HMAC_REG_HMAC384_BLOCK_22                                                                   (32'hd8)
`define CLP_HMAC_REG_HMAC384_BLOCK_23                                                               (32'h100100dc)
`define HMAC_REG_HMAC384_BLOCK_23                                                                   (32'hdc)
`define CLP_HMAC_REG_HMAC384_BLOCK_24                                                               (32'h100100e0)
`define HMAC_REG_HMAC384_BLOCK_24                                                                   (32'he0)
`define CLP_HMAC_REG_HMAC384_BLOCK_25                                                               (32'h100100e4)
`define HMAC_REG_HMAC384_BLOCK_25                                                                   (32'he4)
`define CLP_HMAC_REG_HMAC384_BLOCK_26                                                               (32'h100100e8)
`define HMAC_REG_HMAC384_BLOCK_26                                                                   (32'he8)
`define CLP_HMAC_REG_HMAC384_BLOCK_27                                                               (32'h100100ec)
`define HMAC_REG_HMAC384_BLOCK_27                                                                   (32'hec)
`define CLP_HMAC_REG_HMAC384_BLOCK_28                                                               (32'h100100f0)
`define HMAC_REG_HMAC384_BLOCK_28                                                                   (32'hf0)
`define CLP_HMAC_REG_HMAC384_BLOCK_29                                                               (32'h100100f4)
`define HMAC_REG_HMAC384_BLOCK_29                                                                   (32'hf4)
`define CLP_HMAC_REG_HMAC384_BLOCK_30                                                               (32'h100100f8)
`define HMAC_REG_HMAC384_BLOCK_30                                                                   (32'hf8)
`define CLP_HMAC_REG_HMAC384_BLOCK_31                                                               (32'h100100fc)
`define HMAC_REG_HMAC384_BLOCK_31                                                                   (32'hfc)
`define CLP_HMAC_REG_HMAC384_TAG_0                                                                  (32'h10010100)
`define HMAC_REG_HMAC384_TAG_0                                                                      (32'h100)
`define CLP_HMAC_REG_HMAC384_TAG_1                                                                  (32'h10010104)
`define HMAC_REG_HMAC384_TAG_1                                                                      (32'h104)
`define CLP_HMAC_REG_HMAC384_TAG_2                                                                  (32'h10010108)
`define HMAC_REG_HMAC384_TAG_2                                                                      (32'h108)
`define CLP_HMAC_REG_HMAC384_TAG_3                                                                  (32'h1001010c)
`define HMAC_REG_HMAC384_TAG_3                                                                      (32'h10c)
`define CLP_HMAC_REG_HMAC384_TAG_4                                                                  (32'h10010110)
`define HMAC_REG_HMAC384_TAG_4                                                                      (32'h110)
`define CLP_HMAC_REG_HMAC384_TAG_5                                                                  (32'h10010114)
`define HMAC_REG_HMAC384_TAG_5                                                                      (32'h114)
`define CLP_HMAC_REG_HMAC384_TAG_6                                                                  (32'h10010118)
`define HMAC_REG_HMAC384_TAG_6                                                                      (32'h118)
`define CLP_HMAC_REG_HMAC384_TAG_7                                                                  (32'h1001011c)
`define HMAC_REG_HMAC384_TAG_7                                                                      (32'h11c)
`define CLP_HMAC_REG_HMAC384_TAG_8                                                                  (32'h10010120)
`define HMAC_REG_HMAC384_TAG_8                                                                      (32'h120)
`define CLP_HMAC_REG_HMAC384_TAG_9                                                                  (32'h10010124)
`define HMAC_REG_HMAC384_TAG_9                                                                      (32'h124)
`define CLP_HMAC_REG_HMAC384_TAG_10                                                                 (32'h10010128)
`define HMAC_REG_HMAC384_TAG_10                                                                     (32'h128)
`define CLP_HMAC_REG_HMAC384_TAG_11                                                                 (32'h1001012c)
`define HMAC_REG_HMAC384_TAG_11                                                                     (32'h12c)
`define CLP_HMAC_REG_HMAC384_LFSR_SEED_0                                                            (32'h10010130)
`define HMAC_REG_HMAC384_LFSR_SEED_0                                                                (32'h130)
`define CLP_HMAC_REG_HMAC384_LFSR_SEED_1                                                            (32'h10010134)
`define HMAC_REG_HMAC384_LFSR_SEED_1                                                                (32'h134)
`define CLP_HMAC_REG_HMAC384_LFSR_SEED_2                                                            (32'h10010138)
`define HMAC_REG_HMAC384_LFSR_SEED_2                                                                (32'h138)
`define CLP_HMAC_REG_HMAC384_LFSR_SEED_3                                                            (32'h1001013c)
`define HMAC_REG_HMAC384_LFSR_SEED_3                                                                (32'h13c)
`define CLP_HMAC_REG_HMAC384_LFSR_SEED_4                                                            (32'h10010140)
`define HMAC_REG_HMAC384_LFSR_SEED_4                                                                (32'h140)
`define CLP_HMAC_REG_HMAC384_KV_RD_KEY_CTRL                                                         (32'h10010600)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL                                                             (32'h600)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_READ_EN_LOW                                                 (0)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_READ_EN_MASK                                                (32'h1)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_READ_ENTRY_LOW                                              (1)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_READ_ENTRY_MASK                                             (32'h3e)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_PCR_HASH_EXTEND_LOW                                         (6)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_PCR_HASH_EXTEND_MASK                                        (32'h40)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_RSVD_LOW                                                    (7)
`define HMAC_REG_HMAC384_KV_RD_KEY_CTRL_RSVD_MASK                                                   (32'hffffff80)
`define CLP_HMAC_REG_HMAC384_KV_RD_KEY_STATUS                                                       (32'h10010604)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS                                                           (32'h604)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_READY_LOW                                                 (0)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_READY_MASK                                                (32'h1)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_VALID_LOW                                                 (1)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_VALID_MASK                                                (32'h2)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_ERROR_LOW                                                 (2)
`define HMAC_REG_HMAC384_KV_RD_KEY_STATUS_ERROR_MASK                                                (32'h3fc)
`define CLP_HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL                                                       (32'h10010608)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL                                                           (32'h608)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_READ_EN_LOW                                               (0)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_READ_EN_MASK                                              (32'h1)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_READ_ENTRY_LOW                                            (1)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_READ_ENTRY_MASK                                           (32'h3e)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_PCR_HASH_EXTEND_LOW                                       (6)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_PCR_HASH_EXTEND_MASK                                      (32'h40)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_RSVD_LOW                                                  (7)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_CTRL_RSVD_MASK                                                 (32'hffffff80)
`define CLP_HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS                                                     (32'h1001060c)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS                                                         (32'h60c)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_READY_LOW                                               (0)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_READY_MASK                                              (32'h1)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_VALID_LOW                                               (1)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_VALID_MASK                                              (32'h2)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_ERROR_LOW                                               (2)
`define HMAC_REG_HMAC384_KV_RD_BLOCK_STATUS_ERROR_MASK                                              (32'h3fc)
`define CLP_HMAC_REG_HMAC384_KV_WR_CTRL                                                             (32'h10010610)
`define HMAC_REG_HMAC384_KV_WR_CTRL                                                                 (32'h610)
`define HMAC_REG_HMAC384_KV_WR_CTRL_WRITE_EN_LOW                                                    (0)
`define HMAC_REG_HMAC384_KV_WR_CTRL_WRITE_EN_MASK                                                   (32'h1)
`define HMAC_REG_HMAC384_KV_WR_CTRL_WRITE_ENTRY_LOW                                                 (1)
`define HMAC_REG_HMAC384_KV_WR_CTRL_WRITE_ENTRY_MASK                                                (32'h3e)
`define HMAC_REG_HMAC384_KV_WR_CTRL_HMAC_KEY_DEST_VALID_LOW                                         (6)
`define HMAC_REG_HMAC384_KV_WR_CTRL_HMAC_KEY_DEST_VALID_MASK                                        (32'h40)
`define HMAC_REG_HMAC384_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                       (7)
`define HMAC_REG_HMAC384_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                      (32'h80)
`define HMAC_REG_HMAC384_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_LOW                                        (8)
`define HMAC_REG_HMAC384_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_MASK                                       (32'h100)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_PKEY_DEST_VALID_LOW                                         (9)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_PKEY_DEST_VALID_MASK                                        (32'h200)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_SEED_DEST_VALID_LOW                                         (10)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_SEED_DEST_VALID_MASK                                        (32'h400)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_MSG_DEST_VALID_LOW                                          (11)
`define HMAC_REG_HMAC384_KV_WR_CTRL_ECC_MSG_DEST_VALID_MASK                                         (32'h800)
`define HMAC_REG_HMAC384_KV_WR_CTRL_RSVD_LOW                                                        (12)
`define HMAC_REG_HMAC384_KV_WR_CTRL_RSVD_MASK                                                       (32'hfffff000)
`define CLP_HMAC_REG_HMAC384_KV_WR_STATUS                                                           (32'h10010614)
`define HMAC_REG_HMAC384_KV_WR_STATUS                                                               (32'h614)
`define HMAC_REG_HMAC384_KV_WR_STATUS_READY_LOW                                                     (0)
`define HMAC_REG_HMAC384_KV_WR_STATUS_READY_MASK                                                    (32'h1)
`define HMAC_REG_HMAC384_KV_WR_STATUS_VALID_LOW                                                     (1)
`define HMAC_REG_HMAC384_KV_WR_STATUS_VALID_MASK                                                    (32'h2)
`define HMAC_REG_HMAC384_KV_WR_STATUS_ERROR_LOW                                                     (2)
`define HMAC_REG_HMAC384_KV_WR_STATUS_ERROR_MASK                                                    (32'h3fc)
`define CLP_HMAC_REG_INTR_BLOCK_RF_START                                                            (32'h10010800)
`define CLP_HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                 (32'h10010800)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                     (32'h800)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                        (0)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                       (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                        (1)
`define HMAC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                       (32'h2)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                  (32'h10010804)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                      (32'h804)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                        (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                       (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                        (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                       (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                        (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                       (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                        (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                       (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                  (32'h10010808)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                      (32'h808)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                                (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                               (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                              (32'h1001080c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                  (32'h80c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                      (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                     (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                              (32'h10010810)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                  (32'h810)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                      (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                     (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                            (32'h10010814)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                                (32'h814)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                                 (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                                (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                                 (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                                (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                                 (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                                (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                                 (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                                (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                            (32'h10010818)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                                (32'h818)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                         (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                        (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                (32'h1001081c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                    (32'h81c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                    (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                   (32'h1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                    (1)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                   (32'h2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                    (2)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                   (32'h4)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                    (3)
`define HMAC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                   (32'h8)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                (32'h10010820)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                    (32'h820)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                            (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                           (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                              (32'h10010900)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                  (32'h900)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                              (32'h10010904)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                  (32'h904)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                              (32'h10010908)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                  (32'h908)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                              (32'h1001090c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                  (32'h90c)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                      (32'h10010980)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                          (32'h980)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                         (32'h10010a00)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                             (32'ha00)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                         (32'h10010a04)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                             (32'ha04)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                         (32'h10010a08)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                             (32'ha08)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                         (32'h10010a0c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                             (32'ha0c)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                   (0)
`define HMAC_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                  (32'h1)
`define CLP_HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                 (32'h10010a10)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                     (32'ha10)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                           (0)
`define HMAC_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                          (32'h1)
`define CLP_KV_REG_BASE_ADDR                                                                        (32'h10018000)
`define CLP_KV_REG_KEY_CTRL_0                                                                       (32'h10018000)
`define KV_REG_KEY_CTRL_0                                                                           (32'h0)
`define KV_REG_KEY_CTRL_0_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_0_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_0_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_0_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_0_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_0_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_0_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_0_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_0_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_0_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_0_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_0_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_0_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_0_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_1                                                                       (32'h10018004)
`define KV_REG_KEY_CTRL_1                                                                           (32'h4)
`define KV_REG_KEY_CTRL_1_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_1_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_1_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_1_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_1_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_1_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_1_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_1_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_1_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_1_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_1_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_1_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_1_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_1_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_2                                                                       (32'h10018008)
`define KV_REG_KEY_CTRL_2                                                                           (32'h8)
`define KV_REG_KEY_CTRL_2_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_2_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_2_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_2_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_2_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_2_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_2_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_2_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_2_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_2_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_2_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_2_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_2_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_2_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_3                                                                       (32'h1001800c)
`define KV_REG_KEY_CTRL_3                                                                           (32'hc)
`define KV_REG_KEY_CTRL_3_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_3_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_3_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_3_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_3_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_3_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_3_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_3_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_3_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_3_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_3_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_3_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_3_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_3_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_4                                                                       (32'h10018010)
`define KV_REG_KEY_CTRL_4                                                                           (32'h10)
`define KV_REG_KEY_CTRL_4_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_4_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_4_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_4_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_4_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_4_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_4_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_4_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_4_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_4_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_4_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_4_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_4_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_4_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_5                                                                       (32'h10018014)
`define KV_REG_KEY_CTRL_5                                                                           (32'h14)
`define KV_REG_KEY_CTRL_5_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_5_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_5_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_5_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_5_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_5_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_5_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_5_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_5_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_5_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_5_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_5_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_5_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_5_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_6                                                                       (32'h10018018)
`define KV_REG_KEY_CTRL_6                                                                           (32'h18)
`define KV_REG_KEY_CTRL_6_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_6_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_6_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_6_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_6_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_6_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_6_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_6_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_6_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_6_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_6_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_6_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_6_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_6_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_7                                                                       (32'h1001801c)
`define KV_REG_KEY_CTRL_7                                                                           (32'h1c)
`define KV_REG_KEY_CTRL_7_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_7_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_7_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_7_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_7_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_7_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_7_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_7_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_7_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_7_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_7_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_7_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_7_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_7_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_8                                                                       (32'h10018020)
`define KV_REG_KEY_CTRL_8                                                                           (32'h20)
`define KV_REG_KEY_CTRL_8_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_8_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_8_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_8_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_8_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_8_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_8_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_8_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_8_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_8_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_8_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_8_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_8_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_8_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_9                                                                       (32'h10018024)
`define KV_REG_KEY_CTRL_9                                                                           (32'h24)
`define KV_REG_KEY_CTRL_9_LOCK_WR_LOW                                                               (0)
`define KV_REG_KEY_CTRL_9_LOCK_WR_MASK                                                              (32'h1)
`define KV_REG_KEY_CTRL_9_LOCK_USE_LOW                                                              (1)
`define KV_REG_KEY_CTRL_9_LOCK_USE_MASK                                                             (32'h2)
`define KV_REG_KEY_CTRL_9_CLEAR_LOW                                                                 (2)
`define KV_REG_KEY_CTRL_9_CLEAR_MASK                                                                (32'h4)
`define KV_REG_KEY_CTRL_9_RSVD0_LOW                                                                 (3)
`define KV_REG_KEY_CTRL_9_RSVD0_MASK                                                                (32'h8)
`define KV_REG_KEY_CTRL_9_RSVD1_LOW                                                                 (4)
`define KV_REG_KEY_CTRL_9_RSVD1_MASK                                                                (32'h1f0)
`define KV_REG_KEY_CTRL_9_DEST_VALID_LOW                                                            (9)
`define KV_REG_KEY_CTRL_9_DEST_VALID_MASK                                                           (32'h7e00)
`define KV_REG_KEY_CTRL_9_LAST_DWORD_LOW                                                            (15)
`define KV_REG_KEY_CTRL_9_LAST_DWORD_MASK                                                           (32'h78000)
`define CLP_KV_REG_KEY_CTRL_10                                                                      (32'h10018028)
`define KV_REG_KEY_CTRL_10                                                                          (32'h28)
`define KV_REG_KEY_CTRL_10_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_10_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_10_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_10_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_10_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_10_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_10_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_10_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_10_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_10_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_10_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_10_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_10_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_10_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_11                                                                      (32'h1001802c)
`define KV_REG_KEY_CTRL_11                                                                          (32'h2c)
`define KV_REG_KEY_CTRL_11_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_11_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_11_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_11_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_11_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_11_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_11_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_11_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_11_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_11_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_11_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_11_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_11_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_11_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_12                                                                      (32'h10018030)
`define KV_REG_KEY_CTRL_12                                                                          (32'h30)
`define KV_REG_KEY_CTRL_12_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_12_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_12_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_12_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_12_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_12_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_12_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_12_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_12_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_12_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_12_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_12_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_12_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_12_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_13                                                                      (32'h10018034)
`define KV_REG_KEY_CTRL_13                                                                          (32'h34)
`define KV_REG_KEY_CTRL_13_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_13_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_13_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_13_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_13_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_13_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_13_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_13_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_13_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_13_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_13_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_13_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_13_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_13_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_14                                                                      (32'h10018038)
`define KV_REG_KEY_CTRL_14                                                                          (32'h38)
`define KV_REG_KEY_CTRL_14_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_14_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_14_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_14_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_14_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_14_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_14_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_14_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_14_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_14_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_14_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_14_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_14_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_14_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_15                                                                      (32'h1001803c)
`define KV_REG_KEY_CTRL_15                                                                          (32'h3c)
`define KV_REG_KEY_CTRL_15_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_15_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_15_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_15_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_15_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_15_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_15_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_15_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_15_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_15_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_15_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_15_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_15_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_15_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_16                                                                      (32'h10018040)
`define KV_REG_KEY_CTRL_16                                                                          (32'h40)
`define KV_REG_KEY_CTRL_16_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_16_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_16_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_16_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_16_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_16_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_16_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_16_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_16_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_16_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_16_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_16_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_16_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_16_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_17                                                                      (32'h10018044)
`define KV_REG_KEY_CTRL_17                                                                          (32'h44)
`define KV_REG_KEY_CTRL_17_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_17_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_17_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_17_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_17_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_17_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_17_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_17_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_17_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_17_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_17_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_17_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_17_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_17_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_18                                                                      (32'h10018048)
`define KV_REG_KEY_CTRL_18                                                                          (32'h48)
`define KV_REG_KEY_CTRL_18_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_18_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_18_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_18_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_18_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_18_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_18_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_18_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_18_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_18_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_18_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_18_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_18_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_18_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_19                                                                      (32'h1001804c)
`define KV_REG_KEY_CTRL_19                                                                          (32'h4c)
`define KV_REG_KEY_CTRL_19_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_19_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_19_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_19_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_19_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_19_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_19_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_19_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_19_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_19_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_19_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_19_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_19_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_19_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_20                                                                      (32'h10018050)
`define KV_REG_KEY_CTRL_20                                                                          (32'h50)
`define KV_REG_KEY_CTRL_20_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_20_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_20_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_20_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_20_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_20_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_20_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_20_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_20_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_20_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_20_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_20_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_20_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_20_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_21                                                                      (32'h10018054)
`define KV_REG_KEY_CTRL_21                                                                          (32'h54)
`define KV_REG_KEY_CTRL_21_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_21_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_21_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_21_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_21_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_21_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_21_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_21_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_21_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_21_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_21_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_21_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_21_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_21_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_22                                                                      (32'h10018058)
`define KV_REG_KEY_CTRL_22                                                                          (32'h58)
`define KV_REG_KEY_CTRL_22_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_22_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_22_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_22_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_22_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_22_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_22_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_22_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_22_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_22_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_22_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_22_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_22_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_22_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_23                                                                      (32'h1001805c)
`define KV_REG_KEY_CTRL_23                                                                          (32'h5c)
`define KV_REG_KEY_CTRL_23_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_23_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_23_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_23_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_23_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_23_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_23_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_23_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_23_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_23_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_23_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_23_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_23_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_23_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_24                                                                      (32'h10018060)
`define KV_REG_KEY_CTRL_24                                                                          (32'h60)
`define KV_REG_KEY_CTRL_24_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_24_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_24_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_24_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_24_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_24_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_24_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_24_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_24_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_24_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_24_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_24_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_24_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_24_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_25                                                                      (32'h10018064)
`define KV_REG_KEY_CTRL_25                                                                          (32'h64)
`define KV_REG_KEY_CTRL_25_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_25_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_25_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_25_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_25_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_25_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_25_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_25_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_25_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_25_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_25_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_25_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_25_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_25_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_26                                                                      (32'h10018068)
`define KV_REG_KEY_CTRL_26                                                                          (32'h68)
`define KV_REG_KEY_CTRL_26_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_26_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_26_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_26_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_26_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_26_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_26_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_26_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_26_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_26_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_26_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_26_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_26_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_26_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_27                                                                      (32'h1001806c)
`define KV_REG_KEY_CTRL_27                                                                          (32'h6c)
`define KV_REG_KEY_CTRL_27_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_27_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_27_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_27_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_27_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_27_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_27_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_27_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_27_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_27_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_27_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_27_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_27_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_27_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_28                                                                      (32'h10018070)
`define KV_REG_KEY_CTRL_28                                                                          (32'h70)
`define KV_REG_KEY_CTRL_28_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_28_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_28_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_28_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_28_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_28_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_28_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_28_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_28_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_28_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_28_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_28_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_28_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_28_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_29                                                                      (32'h10018074)
`define KV_REG_KEY_CTRL_29                                                                          (32'h74)
`define KV_REG_KEY_CTRL_29_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_29_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_29_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_29_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_29_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_29_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_29_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_29_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_29_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_29_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_29_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_29_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_29_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_29_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_30                                                                      (32'h10018078)
`define KV_REG_KEY_CTRL_30                                                                          (32'h78)
`define KV_REG_KEY_CTRL_30_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_30_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_30_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_30_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_30_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_30_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_30_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_30_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_30_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_30_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_30_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_30_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_30_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_30_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_CTRL_31                                                                      (32'h1001807c)
`define KV_REG_KEY_CTRL_31                                                                          (32'h7c)
`define KV_REG_KEY_CTRL_31_LOCK_WR_LOW                                                              (0)
`define KV_REG_KEY_CTRL_31_LOCK_WR_MASK                                                             (32'h1)
`define KV_REG_KEY_CTRL_31_LOCK_USE_LOW                                                             (1)
`define KV_REG_KEY_CTRL_31_LOCK_USE_MASK                                                            (32'h2)
`define KV_REG_KEY_CTRL_31_CLEAR_LOW                                                                (2)
`define KV_REG_KEY_CTRL_31_CLEAR_MASK                                                               (32'h4)
`define KV_REG_KEY_CTRL_31_RSVD0_LOW                                                                (3)
`define KV_REG_KEY_CTRL_31_RSVD0_MASK                                                               (32'h8)
`define KV_REG_KEY_CTRL_31_RSVD1_LOW                                                                (4)
`define KV_REG_KEY_CTRL_31_RSVD1_MASK                                                               (32'h1f0)
`define KV_REG_KEY_CTRL_31_DEST_VALID_LOW                                                           (9)
`define KV_REG_KEY_CTRL_31_DEST_VALID_MASK                                                          (32'h7e00)
`define KV_REG_KEY_CTRL_31_LAST_DWORD_LOW                                                           (15)
`define KV_REG_KEY_CTRL_31_LAST_DWORD_MASK                                                          (32'h78000)
`define CLP_KV_REG_KEY_ENTRY_0_0                                                                    (32'h10018600)
`define KV_REG_KEY_ENTRY_0_0                                                                        (32'h600)
`define CLP_KV_REG_KEY_ENTRY_0_1                                                                    (32'h10018604)
`define KV_REG_KEY_ENTRY_0_1                                                                        (32'h604)
`define CLP_KV_REG_KEY_ENTRY_0_2                                                                    (32'h10018608)
`define KV_REG_KEY_ENTRY_0_2                                                                        (32'h608)
`define CLP_KV_REG_KEY_ENTRY_0_3                                                                    (32'h1001860c)
`define KV_REG_KEY_ENTRY_0_3                                                                        (32'h60c)
`define CLP_KV_REG_KEY_ENTRY_0_4                                                                    (32'h10018610)
`define KV_REG_KEY_ENTRY_0_4                                                                        (32'h610)
`define CLP_KV_REG_KEY_ENTRY_0_5                                                                    (32'h10018614)
`define KV_REG_KEY_ENTRY_0_5                                                                        (32'h614)
`define CLP_KV_REG_KEY_ENTRY_0_6                                                                    (32'h10018618)
`define KV_REG_KEY_ENTRY_0_6                                                                        (32'h618)
`define CLP_KV_REG_KEY_ENTRY_0_7                                                                    (32'h1001861c)
`define KV_REG_KEY_ENTRY_0_7                                                                        (32'h61c)
`define CLP_KV_REG_KEY_ENTRY_0_8                                                                    (32'h10018620)
`define KV_REG_KEY_ENTRY_0_8                                                                        (32'h620)
`define CLP_KV_REG_KEY_ENTRY_0_9                                                                    (32'h10018624)
`define KV_REG_KEY_ENTRY_0_9                                                                        (32'h624)
`define CLP_KV_REG_KEY_ENTRY_0_10                                                                   (32'h10018628)
`define KV_REG_KEY_ENTRY_0_10                                                                       (32'h628)
`define CLP_KV_REG_KEY_ENTRY_0_11                                                                   (32'h1001862c)
`define KV_REG_KEY_ENTRY_0_11                                                                       (32'h62c)
`define CLP_KV_REG_KEY_ENTRY_1_0                                                                    (32'h10018630)
`define KV_REG_KEY_ENTRY_1_0                                                                        (32'h630)
`define CLP_KV_REG_KEY_ENTRY_1_1                                                                    (32'h10018634)
`define KV_REG_KEY_ENTRY_1_1                                                                        (32'h634)
`define CLP_KV_REG_KEY_ENTRY_1_2                                                                    (32'h10018638)
`define KV_REG_KEY_ENTRY_1_2                                                                        (32'h638)
`define CLP_KV_REG_KEY_ENTRY_1_3                                                                    (32'h1001863c)
`define KV_REG_KEY_ENTRY_1_3                                                                        (32'h63c)
`define CLP_KV_REG_KEY_ENTRY_1_4                                                                    (32'h10018640)
`define KV_REG_KEY_ENTRY_1_4                                                                        (32'h640)
`define CLP_KV_REG_KEY_ENTRY_1_5                                                                    (32'h10018644)
`define KV_REG_KEY_ENTRY_1_5                                                                        (32'h644)
`define CLP_KV_REG_KEY_ENTRY_1_6                                                                    (32'h10018648)
`define KV_REG_KEY_ENTRY_1_6                                                                        (32'h648)
`define CLP_KV_REG_KEY_ENTRY_1_7                                                                    (32'h1001864c)
`define KV_REG_KEY_ENTRY_1_7                                                                        (32'h64c)
`define CLP_KV_REG_KEY_ENTRY_1_8                                                                    (32'h10018650)
`define KV_REG_KEY_ENTRY_1_8                                                                        (32'h650)
`define CLP_KV_REG_KEY_ENTRY_1_9                                                                    (32'h10018654)
`define KV_REG_KEY_ENTRY_1_9                                                                        (32'h654)
`define CLP_KV_REG_KEY_ENTRY_1_10                                                                   (32'h10018658)
`define KV_REG_KEY_ENTRY_1_10                                                                       (32'h658)
`define CLP_KV_REG_KEY_ENTRY_1_11                                                                   (32'h1001865c)
`define KV_REG_KEY_ENTRY_1_11                                                                       (32'h65c)
`define CLP_KV_REG_KEY_ENTRY_2_0                                                                    (32'h10018660)
`define KV_REG_KEY_ENTRY_2_0                                                                        (32'h660)
`define CLP_KV_REG_KEY_ENTRY_2_1                                                                    (32'h10018664)
`define KV_REG_KEY_ENTRY_2_1                                                                        (32'h664)
`define CLP_KV_REG_KEY_ENTRY_2_2                                                                    (32'h10018668)
`define KV_REG_KEY_ENTRY_2_2                                                                        (32'h668)
`define CLP_KV_REG_KEY_ENTRY_2_3                                                                    (32'h1001866c)
`define KV_REG_KEY_ENTRY_2_3                                                                        (32'h66c)
`define CLP_KV_REG_KEY_ENTRY_2_4                                                                    (32'h10018670)
`define KV_REG_KEY_ENTRY_2_4                                                                        (32'h670)
`define CLP_KV_REG_KEY_ENTRY_2_5                                                                    (32'h10018674)
`define KV_REG_KEY_ENTRY_2_5                                                                        (32'h674)
`define CLP_KV_REG_KEY_ENTRY_2_6                                                                    (32'h10018678)
`define KV_REG_KEY_ENTRY_2_6                                                                        (32'h678)
`define CLP_KV_REG_KEY_ENTRY_2_7                                                                    (32'h1001867c)
`define KV_REG_KEY_ENTRY_2_7                                                                        (32'h67c)
`define CLP_KV_REG_KEY_ENTRY_2_8                                                                    (32'h10018680)
`define KV_REG_KEY_ENTRY_2_8                                                                        (32'h680)
`define CLP_KV_REG_KEY_ENTRY_2_9                                                                    (32'h10018684)
`define KV_REG_KEY_ENTRY_2_9                                                                        (32'h684)
`define CLP_KV_REG_KEY_ENTRY_2_10                                                                   (32'h10018688)
`define KV_REG_KEY_ENTRY_2_10                                                                       (32'h688)
`define CLP_KV_REG_KEY_ENTRY_2_11                                                                   (32'h1001868c)
`define KV_REG_KEY_ENTRY_2_11                                                                       (32'h68c)
`define CLP_KV_REG_KEY_ENTRY_3_0                                                                    (32'h10018690)
`define KV_REG_KEY_ENTRY_3_0                                                                        (32'h690)
`define CLP_KV_REG_KEY_ENTRY_3_1                                                                    (32'h10018694)
`define KV_REG_KEY_ENTRY_3_1                                                                        (32'h694)
`define CLP_KV_REG_KEY_ENTRY_3_2                                                                    (32'h10018698)
`define KV_REG_KEY_ENTRY_3_2                                                                        (32'h698)
`define CLP_KV_REG_KEY_ENTRY_3_3                                                                    (32'h1001869c)
`define KV_REG_KEY_ENTRY_3_3                                                                        (32'h69c)
`define CLP_KV_REG_KEY_ENTRY_3_4                                                                    (32'h100186a0)
`define KV_REG_KEY_ENTRY_3_4                                                                        (32'h6a0)
`define CLP_KV_REG_KEY_ENTRY_3_5                                                                    (32'h100186a4)
`define KV_REG_KEY_ENTRY_3_5                                                                        (32'h6a4)
`define CLP_KV_REG_KEY_ENTRY_3_6                                                                    (32'h100186a8)
`define KV_REG_KEY_ENTRY_3_6                                                                        (32'h6a8)
`define CLP_KV_REG_KEY_ENTRY_3_7                                                                    (32'h100186ac)
`define KV_REG_KEY_ENTRY_3_7                                                                        (32'h6ac)
`define CLP_KV_REG_KEY_ENTRY_3_8                                                                    (32'h100186b0)
`define KV_REG_KEY_ENTRY_3_8                                                                        (32'h6b0)
`define CLP_KV_REG_KEY_ENTRY_3_9                                                                    (32'h100186b4)
`define KV_REG_KEY_ENTRY_3_9                                                                        (32'h6b4)
`define CLP_KV_REG_KEY_ENTRY_3_10                                                                   (32'h100186b8)
`define KV_REG_KEY_ENTRY_3_10                                                                       (32'h6b8)
`define CLP_KV_REG_KEY_ENTRY_3_11                                                                   (32'h100186bc)
`define KV_REG_KEY_ENTRY_3_11                                                                       (32'h6bc)
`define CLP_KV_REG_KEY_ENTRY_4_0                                                                    (32'h100186c0)
`define KV_REG_KEY_ENTRY_4_0                                                                        (32'h6c0)
`define CLP_KV_REG_KEY_ENTRY_4_1                                                                    (32'h100186c4)
`define KV_REG_KEY_ENTRY_4_1                                                                        (32'h6c4)
`define CLP_KV_REG_KEY_ENTRY_4_2                                                                    (32'h100186c8)
`define KV_REG_KEY_ENTRY_4_2                                                                        (32'h6c8)
`define CLP_KV_REG_KEY_ENTRY_4_3                                                                    (32'h100186cc)
`define KV_REG_KEY_ENTRY_4_3                                                                        (32'h6cc)
`define CLP_KV_REG_KEY_ENTRY_4_4                                                                    (32'h100186d0)
`define KV_REG_KEY_ENTRY_4_4                                                                        (32'h6d0)
`define CLP_KV_REG_KEY_ENTRY_4_5                                                                    (32'h100186d4)
`define KV_REG_KEY_ENTRY_4_5                                                                        (32'h6d4)
`define CLP_KV_REG_KEY_ENTRY_4_6                                                                    (32'h100186d8)
`define KV_REG_KEY_ENTRY_4_6                                                                        (32'h6d8)
`define CLP_KV_REG_KEY_ENTRY_4_7                                                                    (32'h100186dc)
`define KV_REG_KEY_ENTRY_4_7                                                                        (32'h6dc)
`define CLP_KV_REG_KEY_ENTRY_4_8                                                                    (32'h100186e0)
`define KV_REG_KEY_ENTRY_4_8                                                                        (32'h6e0)
`define CLP_KV_REG_KEY_ENTRY_4_9                                                                    (32'h100186e4)
`define KV_REG_KEY_ENTRY_4_9                                                                        (32'h6e4)
`define CLP_KV_REG_KEY_ENTRY_4_10                                                                   (32'h100186e8)
`define KV_REG_KEY_ENTRY_4_10                                                                       (32'h6e8)
`define CLP_KV_REG_KEY_ENTRY_4_11                                                                   (32'h100186ec)
`define KV_REG_KEY_ENTRY_4_11                                                                       (32'h6ec)
`define CLP_KV_REG_KEY_ENTRY_5_0                                                                    (32'h100186f0)
`define KV_REG_KEY_ENTRY_5_0                                                                        (32'h6f0)
`define CLP_KV_REG_KEY_ENTRY_5_1                                                                    (32'h100186f4)
`define KV_REG_KEY_ENTRY_5_1                                                                        (32'h6f4)
`define CLP_KV_REG_KEY_ENTRY_5_2                                                                    (32'h100186f8)
`define KV_REG_KEY_ENTRY_5_2                                                                        (32'h6f8)
`define CLP_KV_REG_KEY_ENTRY_5_3                                                                    (32'h100186fc)
`define KV_REG_KEY_ENTRY_5_3                                                                        (32'h6fc)
`define CLP_KV_REG_KEY_ENTRY_5_4                                                                    (32'h10018700)
`define KV_REG_KEY_ENTRY_5_4                                                                        (32'h700)
`define CLP_KV_REG_KEY_ENTRY_5_5                                                                    (32'h10018704)
`define KV_REG_KEY_ENTRY_5_5                                                                        (32'h704)
`define CLP_KV_REG_KEY_ENTRY_5_6                                                                    (32'h10018708)
`define KV_REG_KEY_ENTRY_5_6                                                                        (32'h708)
`define CLP_KV_REG_KEY_ENTRY_5_7                                                                    (32'h1001870c)
`define KV_REG_KEY_ENTRY_5_7                                                                        (32'h70c)
`define CLP_KV_REG_KEY_ENTRY_5_8                                                                    (32'h10018710)
`define KV_REG_KEY_ENTRY_5_8                                                                        (32'h710)
`define CLP_KV_REG_KEY_ENTRY_5_9                                                                    (32'h10018714)
`define KV_REG_KEY_ENTRY_5_9                                                                        (32'h714)
`define CLP_KV_REG_KEY_ENTRY_5_10                                                                   (32'h10018718)
`define KV_REG_KEY_ENTRY_5_10                                                                       (32'h718)
`define CLP_KV_REG_KEY_ENTRY_5_11                                                                   (32'h1001871c)
`define KV_REG_KEY_ENTRY_5_11                                                                       (32'h71c)
`define CLP_KV_REG_KEY_ENTRY_6_0                                                                    (32'h10018720)
`define KV_REG_KEY_ENTRY_6_0                                                                        (32'h720)
`define CLP_KV_REG_KEY_ENTRY_6_1                                                                    (32'h10018724)
`define KV_REG_KEY_ENTRY_6_1                                                                        (32'h724)
`define CLP_KV_REG_KEY_ENTRY_6_2                                                                    (32'h10018728)
`define KV_REG_KEY_ENTRY_6_2                                                                        (32'h728)
`define CLP_KV_REG_KEY_ENTRY_6_3                                                                    (32'h1001872c)
`define KV_REG_KEY_ENTRY_6_3                                                                        (32'h72c)
`define CLP_KV_REG_KEY_ENTRY_6_4                                                                    (32'h10018730)
`define KV_REG_KEY_ENTRY_6_4                                                                        (32'h730)
`define CLP_KV_REG_KEY_ENTRY_6_5                                                                    (32'h10018734)
`define KV_REG_KEY_ENTRY_6_5                                                                        (32'h734)
`define CLP_KV_REG_KEY_ENTRY_6_6                                                                    (32'h10018738)
`define KV_REG_KEY_ENTRY_6_6                                                                        (32'h738)
`define CLP_KV_REG_KEY_ENTRY_6_7                                                                    (32'h1001873c)
`define KV_REG_KEY_ENTRY_6_7                                                                        (32'h73c)
`define CLP_KV_REG_KEY_ENTRY_6_8                                                                    (32'h10018740)
`define KV_REG_KEY_ENTRY_6_8                                                                        (32'h740)
`define CLP_KV_REG_KEY_ENTRY_6_9                                                                    (32'h10018744)
`define KV_REG_KEY_ENTRY_6_9                                                                        (32'h744)
`define CLP_KV_REG_KEY_ENTRY_6_10                                                                   (32'h10018748)
`define KV_REG_KEY_ENTRY_6_10                                                                       (32'h748)
`define CLP_KV_REG_KEY_ENTRY_6_11                                                                   (32'h1001874c)
`define KV_REG_KEY_ENTRY_6_11                                                                       (32'h74c)
`define CLP_KV_REG_KEY_ENTRY_7_0                                                                    (32'h10018750)
`define KV_REG_KEY_ENTRY_7_0                                                                        (32'h750)
`define CLP_KV_REG_KEY_ENTRY_7_1                                                                    (32'h10018754)
`define KV_REG_KEY_ENTRY_7_1                                                                        (32'h754)
`define CLP_KV_REG_KEY_ENTRY_7_2                                                                    (32'h10018758)
`define KV_REG_KEY_ENTRY_7_2                                                                        (32'h758)
`define CLP_KV_REG_KEY_ENTRY_7_3                                                                    (32'h1001875c)
`define KV_REG_KEY_ENTRY_7_3                                                                        (32'h75c)
`define CLP_KV_REG_KEY_ENTRY_7_4                                                                    (32'h10018760)
`define KV_REG_KEY_ENTRY_7_4                                                                        (32'h760)
`define CLP_KV_REG_KEY_ENTRY_7_5                                                                    (32'h10018764)
`define KV_REG_KEY_ENTRY_7_5                                                                        (32'h764)
`define CLP_KV_REG_KEY_ENTRY_7_6                                                                    (32'h10018768)
`define KV_REG_KEY_ENTRY_7_6                                                                        (32'h768)
`define CLP_KV_REG_KEY_ENTRY_7_7                                                                    (32'h1001876c)
`define KV_REG_KEY_ENTRY_7_7                                                                        (32'h76c)
`define CLP_KV_REG_KEY_ENTRY_7_8                                                                    (32'h10018770)
`define KV_REG_KEY_ENTRY_7_8                                                                        (32'h770)
`define CLP_KV_REG_KEY_ENTRY_7_9                                                                    (32'h10018774)
`define KV_REG_KEY_ENTRY_7_9                                                                        (32'h774)
`define CLP_KV_REG_KEY_ENTRY_7_10                                                                   (32'h10018778)
`define KV_REG_KEY_ENTRY_7_10                                                                       (32'h778)
`define CLP_KV_REG_KEY_ENTRY_7_11                                                                   (32'h1001877c)
`define KV_REG_KEY_ENTRY_7_11                                                                       (32'h77c)
`define CLP_KV_REG_KEY_ENTRY_8_0                                                                    (32'h10018780)
`define KV_REG_KEY_ENTRY_8_0                                                                        (32'h780)
`define CLP_KV_REG_KEY_ENTRY_8_1                                                                    (32'h10018784)
`define KV_REG_KEY_ENTRY_8_1                                                                        (32'h784)
`define CLP_KV_REG_KEY_ENTRY_8_2                                                                    (32'h10018788)
`define KV_REG_KEY_ENTRY_8_2                                                                        (32'h788)
`define CLP_KV_REG_KEY_ENTRY_8_3                                                                    (32'h1001878c)
`define KV_REG_KEY_ENTRY_8_3                                                                        (32'h78c)
`define CLP_KV_REG_KEY_ENTRY_8_4                                                                    (32'h10018790)
`define KV_REG_KEY_ENTRY_8_4                                                                        (32'h790)
`define CLP_KV_REG_KEY_ENTRY_8_5                                                                    (32'h10018794)
`define KV_REG_KEY_ENTRY_8_5                                                                        (32'h794)
`define CLP_KV_REG_KEY_ENTRY_8_6                                                                    (32'h10018798)
`define KV_REG_KEY_ENTRY_8_6                                                                        (32'h798)
`define CLP_KV_REG_KEY_ENTRY_8_7                                                                    (32'h1001879c)
`define KV_REG_KEY_ENTRY_8_7                                                                        (32'h79c)
`define CLP_KV_REG_KEY_ENTRY_8_8                                                                    (32'h100187a0)
`define KV_REG_KEY_ENTRY_8_8                                                                        (32'h7a0)
`define CLP_KV_REG_KEY_ENTRY_8_9                                                                    (32'h100187a4)
`define KV_REG_KEY_ENTRY_8_9                                                                        (32'h7a4)
`define CLP_KV_REG_KEY_ENTRY_8_10                                                                   (32'h100187a8)
`define KV_REG_KEY_ENTRY_8_10                                                                       (32'h7a8)
`define CLP_KV_REG_KEY_ENTRY_8_11                                                                   (32'h100187ac)
`define KV_REG_KEY_ENTRY_8_11                                                                       (32'h7ac)
`define CLP_KV_REG_KEY_ENTRY_9_0                                                                    (32'h100187b0)
`define KV_REG_KEY_ENTRY_9_0                                                                        (32'h7b0)
`define CLP_KV_REG_KEY_ENTRY_9_1                                                                    (32'h100187b4)
`define KV_REG_KEY_ENTRY_9_1                                                                        (32'h7b4)
`define CLP_KV_REG_KEY_ENTRY_9_2                                                                    (32'h100187b8)
`define KV_REG_KEY_ENTRY_9_2                                                                        (32'h7b8)
`define CLP_KV_REG_KEY_ENTRY_9_3                                                                    (32'h100187bc)
`define KV_REG_KEY_ENTRY_9_3                                                                        (32'h7bc)
`define CLP_KV_REG_KEY_ENTRY_9_4                                                                    (32'h100187c0)
`define KV_REG_KEY_ENTRY_9_4                                                                        (32'h7c0)
`define CLP_KV_REG_KEY_ENTRY_9_5                                                                    (32'h100187c4)
`define KV_REG_KEY_ENTRY_9_5                                                                        (32'h7c4)
`define CLP_KV_REG_KEY_ENTRY_9_6                                                                    (32'h100187c8)
`define KV_REG_KEY_ENTRY_9_6                                                                        (32'h7c8)
`define CLP_KV_REG_KEY_ENTRY_9_7                                                                    (32'h100187cc)
`define KV_REG_KEY_ENTRY_9_7                                                                        (32'h7cc)
`define CLP_KV_REG_KEY_ENTRY_9_8                                                                    (32'h100187d0)
`define KV_REG_KEY_ENTRY_9_8                                                                        (32'h7d0)
`define CLP_KV_REG_KEY_ENTRY_9_9                                                                    (32'h100187d4)
`define KV_REG_KEY_ENTRY_9_9                                                                        (32'h7d4)
`define CLP_KV_REG_KEY_ENTRY_9_10                                                                   (32'h100187d8)
`define KV_REG_KEY_ENTRY_9_10                                                                       (32'h7d8)
`define CLP_KV_REG_KEY_ENTRY_9_11                                                                   (32'h100187dc)
`define KV_REG_KEY_ENTRY_9_11                                                                       (32'h7dc)
`define CLP_KV_REG_KEY_ENTRY_10_0                                                                   (32'h100187e0)
`define KV_REG_KEY_ENTRY_10_0                                                                       (32'h7e0)
`define CLP_KV_REG_KEY_ENTRY_10_1                                                                   (32'h100187e4)
`define KV_REG_KEY_ENTRY_10_1                                                                       (32'h7e4)
`define CLP_KV_REG_KEY_ENTRY_10_2                                                                   (32'h100187e8)
`define KV_REG_KEY_ENTRY_10_2                                                                       (32'h7e8)
`define CLP_KV_REG_KEY_ENTRY_10_3                                                                   (32'h100187ec)
`define KV_REG_KEY_ENTRY_10_3                                                                       (32'h7ec)
`define CLP_KV_REG_KEY_ENTRY_10_4                                                                   (32'h100187f0)
`define KV_REG_KEY_ENTRY_10_4                                                                       (32'h7f0)
`define CLP_KV_REG_KEY_ENTRY_10_5                                                                   (32'h100187f4)
`define KV_REG_KEY_ENTRY_10_5                                                                       (32'h7f4)
`define CLP_KV_REG_KEY_ENTRY_10_6                                                                   (32'h100187f8)
`define KV_REG_KEY_ENTRY_10_6                                                                       (32'h7f8)
`define CLP_KV_REG_KEY_ENTRY_10_7                                                                   (32'h100187fc)
`define KV_REG_KEY_ENTRY_10_7                                                                       (32'h7fc)
`define CLP_KV_REG_KEY_ENTRY_10_8                                                                   (32'h10018800)
`define KV_REG_KEY_ENTRY_10_8                                                                       (32'h800)
`define CLP_KV_REG_KEY_ENTRY_10_9                                                                   (32'h10018804)
`define KV_REG_KEY_ENTRY_10_9                                                                       (32'h804)
`define CLP_KV_REG_KEY_ENTRY_10_10                                                                  (32'h10018808)
`define KV_REG_KEY_ENTRY_10_10                                                                      (32'h808)
`define CLP_KV_REG_KEY_ENTRY_10_11                                                                  (32'h1001880c)
`define KV_REG_KEY_ENTRY_10_11                                                                      (32'h80c)
`define CLP_KV_REG_KEY_ENTRY_11_0                                                                   (32'h10018810)
`define KV_REG_KEY_ENTRY_11_0                                                                       (32'h810)
`define CLP_KV_REG_KEY_ENTRY_11_1                                                                   (32'h10018814)
`define KV_REG_KEY_ENTRY_11_1                                                                       (32'h814)
`define CLP_KV_REG_KEY_ENTRY_11_2                                                                   (32'h10018818)
`define KV_REG_KEY_ENTRY_11_2                                                                       (32'h818)
`define CLP_KV_REG_KEY_ENTRY_11_3                                                                   (32'h1001881c)
`define KV_REG_KEY_ENTRY_11_3                                                                       (32'h81c)
`define CLP_KV_REG_KEY_ENTRY_11_4                                                                   (32'h10018820)
`define KV_REG_KEY_ENTRY_11_4                                                                       (32'h820)
`define CLP_KV_REG_KEY_ENTRY_11_5                                                                   (32'h10018824)
`define KV_REG_KEY_ENTRY_11_5                                                                       (32'h824)
`define CLP_KV_REG_KEY_ENTRY_11_6                                                                   (32'h10018828)
`define KV_REG_KEY_ENTRY_11_6                                                                       (32'h828)
`define CLP_KV_REG_KEY_ENTRY_11_7                                                                   (32'h1001882c)
`define KV_REG_KEY_ENTRY_11_7                                                                       (32'h82c)
`define CLP_KV_REG_KEY_ENTRY_11_8                                                                   (32'h10018830)
`define KV_REG_KEY_ENTRY_11_8                                                                       (32'h830)
`define CLP_KV_REG_KEY_ENTRY_11_9                                                                   (32'h10018834)
`define KV_REG_KEY_ENTRY_11_9                                                                       (32'h834)
`define CLP_KV_REG_KEY_ENTRY_11_10                                                                  (32'h10018838)
`define KV_REG_KEY_ENTRY_11_10                                                                      (32'h838)
`define CLP_KV_REG_KEY_ENTRY_11_11                                                                  (32'h1001883c)
`define KV_REG_KEY_ENTRY_11_11                                                                      (32'h83c)
`define CLP_KV_REG_KEY_ENTRY_12_0                                                                   (32'h10018840)
`define KV_REG_KEY_ENTRY_12_0                                                                       (32'h840)
`define CLP_KV_REG_KEY_ENTRY_12_1                                                                   (32'h10018844)
`define KV_REG_KEY_ENTRY_12_1                                                                       (32'h844)
`define CLP_KV_REG_KEY_ENTRY_12_2                                                                   (32'h10018848)
`define KV_REG_KEY_ENTRY_12_2                                                                       (32'h848)
`define CLP_KV_REG_KEY_ENTRY_12_3                                                                   (32'h1001884c)
`define KV_REG_KEY_ENTRY_12_3                                                                       (32'h84c)
`define CLP_KV_REG_KEY_ENTRY_12_4                                                                   (32'h10018850)
`define KV_REG_KEY_ENTRY_12_4                                                                       (32'h850)
`define CLP_KV_REG_KEY_ENTRY_12_5                                                                   (32'h10018854)
`define KV_REG_KEY_ENTRY_12_5                                                                       (32'h854)
`define CLP_KV_REG_KEY_ENTRY_12_6                                                                   (32'h10018858)
`define KV_REG_KEY_ENTRY_12_6                                                                       (32'h858)
`define CLP_KV_REG_KEY_ENTRY_12_7                                                                   (32'h1001885c)
`define KV_REG_KEY_ENTRY_12_7                                                                       (32'h85c)
`define CLP_KV_REG_KEY_ENTRY_12_8                                                                   (32'h10018860)
`define KV_REG_KEY_ENTRY_12_8                                                                       (32'h860)
`define CLP_KV_REG_KEY_ENTRY_12_9                                                                   (32'h10018864)
`define KV_REG_KEY_ENTRY_12_9                                                                       (32'h864)
`define CLP_KV_REG_KEY_ENTRY_12_10                                                                  (32'h10018868)
`define KV_REG_KEY_ENTRY_12_10                                                                      (32'h868)
`define CLP_KV_REG_KEY_ENTRY_12_11                                                                  (32'h1001886c)
`define KV_REG_KEY_ENTRY_12_11                                                                      (32'h86c)
`define CLP_KV_REG_KEY_ENTRY_13_0                                                                   (32'h10018870)
`define KV_REG_KEY_ENTRY_13_0                                                                       (32'h870)
`define CLP_KV_REG_KEY_ENTRY_13_1                                                                   (32'h10018874)
`define KV_REG_KEY_ENTRY_13_1                                                                       (32'h874)
`define CLP_KV_REG_KEY_ENTRY_13_2                                                                   (32'h10018878)
`define KV_REG_KEY_ENTRY_13_2                                                                       (32'h878)
`define CLP_KV_REG_KEY_ENTRY_13_3                                                                   (32'h1001887c)
`define KV_REG_KEY_ENTRY_13_3                                                                       (32'h87c)
`define CLP_KV_REG_KEY_ENTRY_13_4                                                                   (32'h10018880)
`define KV_REG_KEY_ENTRY_13_4                                                                       (32'h880)
`define CLP_KV_REG_KEY_ENTRY_13_5                                                                   (32'h10018884)
`define KV_REG_KEY_ENTRY_13_5                                                                       (32'h884)
`define CLP_KV_REG_KEY_ENTRY_13_6                                                                   (32'h10018888)
`define KV_REG_KEY_ENTRY_13_6                                                                       (32'h888)
`define CLP_KV_REG_KEY_ENTRY_13_7                                                                   (32'h1001888c)
`define KV_REG_KEY_ENTRY_13_7                                                                       (32'h88c)
`define CLP_KV_REG_KEY_ENTRY_13_8                                                                   (32'h10018890)
`define KV_REG_KEY_ENTRY_13_8                                                                       (32'h890)
`define CLP_KV_REG_KEY_ENTRY_13_9                                                                   (32'h10018894)
`define KV_REG_KEY_ENTRY_13_9                                                                       (32'h894)
`define CLP_KV_REG_KEY_ENTRY_13_10                                                                  (32'h10018898)
`define KV_REG_KEY_ENTRY_13_10                                                                      (32'h898)
`define CLP_KV_REG_KEY_ENTRY_13_11                                                                  (32'h1001889c)
`define KV_REG_KEY_ENTRY_13_11                                                                      (32'h89c)
`define CLP_KV_REG_KEY_ENTRY_14_0                                                                   (32'h100188a0)
`define KV_REG_KEY_ENTRY_14_0                                                                       (32'h8a0)
`define CLP_KV_REG_KEY_ENTRY_14_1                                                                   (32'h100188a4)
`define KV_REG_KEY_ENTRY_14_1                                                                       (32'h8a4)
`define CLP_KV_REG_KEY_ENTRY_14_2                                                                   (32'h100188a8)
`define KV_REG_KEY_ENTRY_14_2                                                                       (32'h8a8)
`define CLP_KV_REG_KEY_ENTRY_14_3                                                                   (32'h100188ac)
`define KV_REG_KEY_ENTRY_14_3                                                                       (32'h8ac)
`define CLP_KV_REG_KEY_ENTRY_14_4                                                                   (32'h100188b0)
`define KV_REG_KEY_ENTRY_14_4                                                                       (32'h8b0)
`define CLP_KV_REG_KEY_ENTRY_14_5                                                                   (32'h100188b4)
`define KV_REG_KEY_ENTRY_14_5                                                                       (32'h8b4)
`define CLP_KV_REG_KEY_ENTRY_14_6                                                                   (32'h100188b8)
`define KV_REG_KEY_ENTRY_14_6                                                                       (32'h8b8)
`define CLP_KV_REG_KEY_ENTRY_14_7                                                                   (32'h100188bc)
`define KV_REG_KEY_ENTRY_14_7                                                                       (32'h8bc)
`define CLP_KV_REG_KEY_ENTRY_14_8                                                                   (32'h100188c0)
`define KV_REG_KEY_ENTRY_14_8                                                                       (32'h8c0)
`define CLP_KV_REG_KEY_ENTRY_14_9                                                                   (32'h100188c4)
`define KV_REG_KEY_ENTRY_14_9                                                                       (32'h8c4)
`define CLP_KV_REG_KEY_ENTRY_14_10                                                                  (32'h100188c8)
`define KV_REG_KEY_ENTRY_14_10                                                                      (32'h8c8)
`define CLP_KV_REG_KEY_ENTRY_14_11                                                                  (32'h100188cc)
`define KV_REG_KEY_ENTRY_14_11                                                                      (32'h8cc)
`define CLP_KV_REG_KEY_ENTRY_15_0                                                                   (32'h100188d0)
`define KV_REG_KEY_ENTRY_15_0                                                                       (32'h8d0)
`define CLP_KV_REG_KEY_ENTRY_15_1                                                                   (32'h100188d4)
`define KV_REG_KEY_ENTRY_15_1                                                                       (32'h8d4)
`define CLP_KV_REG_KEY_ENTRY_15_2                                                                   (32'h100188d8)
`define KV_REG_KEY_ENTRY_15_2                                                                       (32'h8d8)
`define CLP_KV_REG_KEY_ENTRY_15_3                                                                   (32'h100188dc)
`define KV_REG_KEY_ENTRY_15_3                                                                       (32'h8dc)
`define CLP_KV_REG_KEY_ENTRY_15_4                                                                   (32'h100188e0)
`define KV_REG_KEY_ENTRY_15_4                                                                       (32'h8e0)
`define CLP_KV_REG_KEY_ENTRY_15_5                                                                   (32'h100188e4)
`define KV_REG_KEY_ENTRY_15_5                                                                       (32'h8e4)
`define CLP_KV_REG_KEY_ENTRY_15_6                                                                   (32'h100188e8)
`define KV_REG_KEY_ENTRY_15_6                                                                       (32'h8e8)
`define CLP_KV_REG_KEY_ENTRY_15_7                                                                   (32'h100188ec)
`define KV_REG_KEY_ENTRY_15_7                                                                       (32'h8ec)
`define CLP_KV_REG_KEY_ENTRY_15_8                                                                   (32'h100188f0)
`define KV_REG_KEY_ENTRY_15_8                                                                       (32'h8f0)
`define CLP_KV_REG_KEY_ENTRY_15_9                                                                   (32'h100188f4)
`define KV_REG_KEY_ENTRY_15_9                                                                       (32'h8f4)
`define CLP_KV_REG_KEY_ENTRY_15_10                                                                  (32'h100188f8)
`define KV_REG_KEY_ENTRY_15_10                                                                      (32'h8f8)
`define CLP_KV_REG_KEY_ENTRY_15_11                                                                  (32'h100188fc)
`define KV_REG_KEY_ENTRY_15_11                                                                      (32'h8fc)
`define CLP_KV_REG_KEY_ENTRY_16_0                                                                   (32'h10018900)
`define KV_REG_KEY_ENTRY_16_0                                                                       (32'h900)
`define CLP_KV_REG_KEY_ENTRY_16_1                                                                   (32'h10018904)
`define KV_REG_KEY_ENTRY_16_1                                                                       (32'h904)
`define CLP_KV_REG_KEY_ENTRY_16_2                                                                   (32'h10018908)
`define KV_REG_KEY_ENTRY_16_2                                                                       (32'h908)
`define CLP_KV_REG_KEY_ENTRY_16_3                                                                   (32'h1001890c)
`define KV_REG_KEY_ENTRY_16_3                                                                       (32'h90c)
`define CLP_KV_REG_KEY_ENTRY_16_4                                                                   (32'h10018910)
`define KV_REG_KEY_ENTRY_16_4                                                                       (32'h910)
`define CLP_KV_REG_KEY_ENTRY_16_5                                                                   (32'h10018914)
`define KV_REG_KEY_ENTRY_16_5                                                                       (32'h914)
`define CLP_KV_REG_KEY_ENTRY_16_6                                                                   (32'h10018918)
`define KV_REG_KEY_ENTRY_16_6                                                                       (32'h918)
`define CLP_KV_REG_KEY_ENTRY_16_7                                                                   (32'h1001891c)
`define KV_REG_KEY_ENTRY_16_7                                                                       (32'h91c)
`define CLP_KV_REG_KEY_ENTRY_16_8                                                                   (32'h10018920)
`define KV_REG_KEY_ENTRY_16_8                                                                       (32'h920)
`define CLP_KV_REG_KEY_ENTRY_16_9                                                                   (32'h10018924)
`define KV_REG_KEY_ENTRY_16_9                                                                       (32'h924)
`define CLP_KV_REG_KEY_ENTRY_16_10                                                                  (32'h10018928)
`define KV_REG_KEY_ENTRY_16_10                                                                      (32'h928)
`define CLP_KV_REG_KEY_ENTRY_16_11                                                                  (32'h1001892c)
`define KV_REG_KEY_ENTRY_16_11                                                                      (32'h92c)
`define CLP_KV_REG_KEY_ENTRY_17_0                                                                   (32'h10018930)
`define KV_REG_KEY_ENTRY_17_0                                                                       (32'h930)
`define CLP_KV_REG_KEY_ENTRY_17_1                                                                   (32'h10018934)
`define KV_REG_KEY_ENTRY_17_1                                                                       (32'h934)
`define CLP_KV_REG_KEY_ENTRY_17_2                                                                   (32'h10018938)
`define KV_REG_KEY_ENTRY_17_2                                                                       (32'h938)
`define CLP_KV_REG_KEY_ENTRY_17_3                                                                   (32'h1001893c)
`define KV_REG_KEY_ENTRY_17_3                                                                       (32'h93c)
`define CLP_KV_REG_KEY_ENTRY_17_4                                                                   (32'h10018940)
`define KV_REG_KEY_ENTRY_17_4                                                                       (32'h940)
`define CLP_KV_REG_KEY_ENTRY_17_5                                                                   (32'h10018944)
`define KV_REG_KEY_ENTRY_17_5                                                                       (32'h944)
`define CLP_KV_REG_KEY_ENTRY_17_6                                                                   (32'h10018948)
`define KV_REG_KEY_ENTRY_17_6                                                                       (32'h948)
`define CLP_KV_REG_KEY_ENTRY_17_7                                                                   (32'h1001894c)
`define KV_REG_KEY_ENTRY_17_7                                                                       (32'h94c)
`define CLP_KV_REG_KEY_ENTRY_17_8                                                                   (32'h10018950)
`define KV_REG_KEY_ENTRY_17_8                                                                       (32'h950)
`define CLP_KV_REG_KEY_ENTRY_17_9                                                                   (32'h10018954)
`define KV_REG_KEY_ENTRY_17_9                                                                       (32'h954)
`define CLP_KV_REG_KEY_ENTRY_17_10                                                                  (32'h10018958)
`define KV_REG_KEY_ENTRY_17_10                                                                      (32'h958)
`define CLP_KV_REG_KEY_ENTRY_17_11                                                                  (32'h1001895c)
`define KV_REG_KEY_ENTRY_17_11                                                                      (32'h95c)
`define CLP_KV_REG_KEY_ENTRY_18_0                                                                   (32'h10018960)
`define KV_REG_KEY_ENTRY_18_0                                                                       (32'h960)
`define CLP_KV_REG_KEY_ENTRY_18_1                                                                   (32'h10018964)
`define KV_REG_KEY_ENTRY_18_1                                                                       (32'h964)
`define CLP_KV_REG_KEY_ENTRY_18_2                                                                   (32'h10018968)
`define KV_REG_KEY_ENTRY_18_2                                                                       (32'h968)
`define CLP_KV_REG_KEY_ENTRY_18_3                                                                   (32'h1001896c)
`define KV_REG_KEY_ENTRY_18_3                                                                       (32'h96c)
`define CLP_KV_REG_KEY_ENTRY_18_4                                                                   (32'h10018970)
`define KV_REG_KEY_ENTRY_18_4                                                                       (32'h970)
`define CLP_KV_REG_KEY_ENTRY_18_5                                                                   (32'h10018974)
`define KV_REG_KEY_ENTRY_18_5                                                                       (32'h974)
`define CLP_KV_REG_KEY_ENTRY_18_6                                                                   (32'h10018978)
`define KV_REG_KEY_ENTRY_18_6                                                                       (32'h978)
`define CLP_KV_REG_KEY_ENTRY_18_7                                                                   (32'h1001897c)
`define KV_REG_KEY_ENTRY_18_7                                                                       (32'h97c)
`define CLP_KV_REG_KEY_ENTRY_18_8                                                                   (32'h10018980)
`define KV_REG_KEY_ENTRY_18_8                                                                       (32'h980)
`define CLP_KV_REG_KEY_ENTRY_18_9                                                                   (32'h10018984)
`define KV_REG_KEY_ENTRY_18_9                                                                       (32'h984)
`define CLP_KV_REG_KEY_ENTRY_18_10                                                                  (32'h10018988)
`define KV_REG_KEY_ENTRY_18_10                                                                      (32'h988)
`define CLP_KV_REG_KEY_ENTRY_18_11                                                                  (32'h1001898c)
`define KV_REG_KEY_ENTRY_18_11                                                                      (32'h98c)
`define CLP_KV_REG_KEY_ENTRY_19_0                                                                   (32'h10018990)
`define KV_REG_KEY_ENTRY_19_0                                                                       (32'h990)
`define CLP_KV_REG_KEY_ENTRY_19_1                                                                   (32'h10018994)
`define KV_REG_KEY_ENTRY_19_1                                                                       (32'h994)
`define CLP_KV_REG_KEY_ENTRY_19_2                                                                   (32'h10018998)
`define KV_REG_KEY_ENTRY_19_2                                                                       (32'h998)
`define CLP_KV_REG_KEY_ENTRY_19_3                                                                   (32'h1001899c)
`define KV_REG_KEY_ENTRY_19_3                                                                       (32'h99c)
`define CLP_KV_REG_KEY_ENTRY_19_4                                                                   (32'h100189a0)
`define KV_REG_KEY_ENTRY_19_4                                                                       (32'h9a0)
`define CLP_KV_REG_KEY_ENTRY_19_5                                                                   (32'h100189a4)
`define KV_REG_KEY_ENTRY_19_5                                                                       (32'h9a4)
`define CLP_KV_REG_KEY_ENTRY_19_6                                                                   (32'h100189a8)
`define KV_REG_KEY_ENTRY_19_6                                                                       (32'h9a8)
`define CLP_KV_REG_KEY_ENTRY_19_7                                                                   (32'h100189ac)
`define KV_REG_KEY_ENTRY_19_7                                                                       (32'h9ac)
`define CLP_KV_REG_KEY_ENTRY_19_8                                                                   (32'h100189b0)
`define KV_REG_KEY_ENTRY_19_8                                                                       (32'h9b0)
`define CLP_KV_REG_KEY_ENTRY_19_9                                                                   (32'h100189b4)
`define KV_REG_KEY_ENTRY_19_9                                                                       (32'h9b4)
`define CLP_KV_REG_KEY_ENTRY_19_10                                                                  (32'h100189b8)
`define KV_REG_KEY_ENTRY_19_10                                                                      (32'h9b8)
`define CLP_KV_REG_KEY_ENTRY_19_11                                                                  (32'h100189bc)
`define KV_REG_KEY_ENTRY_19_11                                                                      (32'h9bc)
`define CLP_KV_REG_KEY_ENTRY_20_0                                                                   (32'h100189c0)
`define KV_REG_KEY_ENTRY_20_0                                                                       (32'h9c0)
`define CLP_KV_REG_KEY_ENTRY_20_1                                                                   (32'h100189c4)
`define KV_REG_KEY_ENTRY_20_1                                                                       (32'h9c4)
`define CLP_KV_REG_KEY_ENTRY_20_2                                                                   (32'h100189c8)
`define KV_REG_KEY_ENTRY_20_2                                                                       (32'h9c8)
`define CLP_KV_REG_KEY_ENTRY_20_3                                                                   (32'h100189cc)
`define KV_REG_KEY_ENTRY_20_3                                                                       (32'h9cc)
`define CLP_KV_REG_KEY_ENTRY_20_4                                                                   (32'h100189d0)
`define KV_REG_KEY_ENTRY_20_4                                                                       (32'h9d0)
`define CLP_KV_REG_KEY_ENTRY_20_5                                                                   (32'h100189d4)
`define KV_REG_KEY_ENTRY_20_5                                                                       (32'h9d4)
`define CLP_KV_REG_KEY_ENTRY_20_6                                                                   (32'h100189d8)
`define KV_REG_KEY_ENTRY_20_6                                                                       (32'h9d8)
`define CLP_KV_REG_KEY_ENTRY_20_7                                                                   (32'h100189dc)
`define KV_REG_KEY_ENTRY_20_7                                                                       (32'h9dc)
`define CLP_KV_REG_KEY_ENTRY_20_8                                                                   (32'h100189e0)
`define KV_REG_KEY_ENTRY_20_8                                                                       (32'h9e0)
`define CLP_KV_REG_KEY_ENTRY_20_9                                                                   (32'h100189e4)
`define KV_REG_KEY_ENTRY_20_9                                                                       (32'h9e4)
`define CLP_KV_REG_KEY_ENTRY_20_10                                                                  (32'h100189e8)
`define KV_REG_KEY_ENTRY_20_10                                                                      (32'h9e8)
`define CLP_KV_REG_KEY_ENTRY_20_11                                                                  (32'h100189ec)
`define KV_REG_KEY_ENTRY_20_11                                                                      (32'h9ec)
`define CLP_KV_REG_KEY_ENTRY_21_0                                                                   (32'h100189f0)
`define KV_REG_KEY_ENTRY_21_0                                                                       (32'h9f0)
`define CLP_KV_REG_KEY_ENTRY_21_1                                                                   (32'h100189f4)
`define KV_REG_KEY_ENTRY_21_1                                                                       (32'h9f4)
`define CLP_KV_REG_KEY_ENTRY_21_2                                                                   (32'h100189f8)
`define KV_REG_KEY_ENTRY_21_2                                                                       (32'h9f8)
`define CLP_KV_REG_KEY_ENTRY_21_3                                                                   (32'h100189fc)
`define KV_REG_KEY_ENTRY_21_3                                                                       (32'h9fc)
`define CLP_KV_REG_KEY_ENTRY_21_4                                                                   (32'h10018a00)
`define KV_REG_KEY_ENTRY_21_4                                                                       (32'ha00)
`define CLP_KV_REG_KEY_ENTRY_21_5                                                                   (32'h10018a04)
`define KV_REG_KEY_ENTRY_21_5                                                                       (32'ha04)
`define CLP_KV_REG_KEY_ENTRY_21_6                                                                   (32'h10018a08)
`define KV_REG_KEY_ENTRY_21_6                                                                       (32'ha08)
`define CLP_KV_REG_KEY_ENTRY_21_7                                                                   (32'h10018a0c)
`define KV_REG_KEY_ENTRY_21_7                                                                       (32'ha0c)
`define CLP_KV_REG_KEY_ENTRY_21_8                                                                   (32'h10018a10)
`define KV_REG_KEY_ENTRY_21_8                                                                       (32'ha10)
`define CLP_KV_REG_KEY_ENTRY_21_9                                                                   (32'h10018a14)
`define KV_REG_KEY_ENTRY_21_9                                                                       (32'ha14)
`define CLP_KV_REG_KEY_ENTRY_21_10                                                                  (32'h10018a18)
`define KV_REG_KEY_ENTRY_21_10                                                                      (32'ha18)
`define CLP_KV_REG_KEY_ENTRY_21_11                                                                  (32'h10018a1c)
`define KV_REG_KEY_ENTRY_21_11                                                                      (32'ha1c)
`define CLP_KV_REG_KEY_ENTRY_22_0                                                                   (32'h10018a20)
`define KV_REG_KEY_ENTRY_22_0                                                                       (32'ha20)
`define CLP_KV_REG_KEY_ENTRY_22_1                                                                   (32'h10018a24)
`define KV_REG_KEY_ENTRY_22_1                                                                       (32'ha24)
`define CLP_KV_REG_KEY_ENTRY_22_2                                                                   (32'h10018a28)
`define KV_REG_KEY_ENTRY_22_2                                                                       (32'ha28)
`define CLP_KV_REG_KEY_ENTRY_22_3                                                                   (32'h10018a2c)
`define KV_REG_KEY_ENTRY_22_3                                                                       (32'ha2c)
`define CLP_KV_REG_KEY_ENTRY_22_4                                                                   (32'h10018a30)
`define KV_REG_KEY_ENTRY_22_4                                                                       (32'ha30)
`define CLP_KV_REG_KEY_ENTRY_22_5                                                                   (32'h10018a34)
`define KV_REG_KEY_ENTRY_22_5                                                                       (32'ha34)
`define CLP_KV_REG_KEY_ENTRY_22_6                                                                   (32'h10018a38)
`define KV_REG_KEY_ENTRY_22_6                                                                       (32'ha38)
`define CLP_KV_REG_KEY_ENTRY_22_7                                                                   (32'h10018a3c)
`define KV_REG_KEY_ENTRY_22_7                                                                       (32'ha3c)
`define CLP_KV_REG_KEY_ENTRY_22_8                                                                   (32'h10018a40)
`define KV_REG_KEY_ENTRY_22_8                                                                       (32'ha40)
`define CLP_KV_REG_KEY_ENTRY_22_9                                                                   (32'h10018a44)
`define KV_REG_KEY_ENTRY_22_9                                                                       (32'ha44)
`define CLP_KV_REG_KEY_ENTRY_22_10                                                                  (32'h10018a48)
`define KV_REG_KEY_ENTRY_22_10                                                                      (32'ha48)
`define CLP_KV_REG_KEY_ENTRY_22_11                                                                  (32'h10018a4c)
`define KV_REG_KEY_ENTRY_22_11                                                                      (32'ha4c)
`define CLP_KV_REG_KEY_ENTRY_23_0                                                                   (32'h10018a50)
`define KV_REG_KEY_ENTRY_23_0                                                                       (32'ha50)
`define CLP_KV_REG_KEY_ENTRY_23_1                                                                   (32'h10018a54)
`define KV_REG_KEY_ENTRY_23_1                                                                       (32'ha54)
`define CLP_KV_REG_KEY_ENTRY_23_2                                                                   (32'h10018a58)
`define KV_REG_KEY_ENTRY_23_2                                                                       (32'ha58)
`define CLP_KV_REG_KEY_ENTRY_23_3                                                                   (32'h10018a5c)
`define KV_REG_KEY_ENTRY_23_3                                                                       (32'ha5c)
`define CLP_KV_REG_KEY_ENTRY_23_4                                                                   (32'h10018a60)
`define KV_REG_KEY_ENTRY_23_4                                                                       (32'ha60)
`define CLP_KV_REG_KEY_ENTRY_23_5                                                                   (32'h10018a64)
`define KV_REG_KEY_ENTRY_23_5                                                                       (32'ha64)
`define CLP_KV_REG_KEY_ENTRY_23_6                                                                   (32'h10018a68)
`define KV_REG_KEY_ENTRY_23_6                                                                       (32'ha68)
`define CLP_KV_REG_KEY_ENTRY_23_7                                                                   (32'h10018a6c)
`define KV_REG_KEY_ENTRY_23_7                                                                       (32'ha6c)
`define CLP_KV_REG_KEY_ENTRY_23_8                                                                   (32'h10018a70)
`define KV_REG_KEY_ENTRY_23_8                                                                       (32'ha70)
`define CLP_KV_REG_KEY_ENTRY_23_9                                                                   (32'h10018a74)
`define KV_REG_KEY_ENTRY_23_9                                                                       (32'ha74)
`define CLP_KV_REG_KEY_ENTRY_23_10                                                                  (32'h10018a78)
`define KV_REG_KEY_ENTRY_23_10                                                                      (32'ha78)
`define CLP_KV_REG_KEY_ENTRY_23_11                                                                  (32'h10018a7c)
`define KV_REG_KEY_ENTRY_23_11                                                                      (32'ha7c)
`define CLP_KV_REG_KEY_ENTRY_24_0                                                                   (32'h10018a80)
`define KV_REG_KEY_ENTRY_24_0                                                                       (32'ha80)
`define CLP_KV_REG_KEY_ENTRY_24_1                                                                   (32'h10018a84)
`define KV_REG_KEY_ENTRY_24_1                                                                       (32'ha84)
`define CLP_KV_REG_KEY_ENTRY_24_2                                                                   (32'h10018a88)
`define KV_REG_KEY_ENTRY_24_2                                                                       (32'ha88)
`define CLP_KV_REG_KEY_ENTRY_24_3                                                                   (32'h10018a8c)
`define KV_REG_KEY_ENTRY_24_3                                                                       (32'ha8c)
`define CLP_KV_REG_KEY_ENTRY_24_4                                                                   (32'h10018a90)
`define KV_REG_KEY_ENTRY_24_4                                                                       (32'ha90)
`define CLP_KV_REG_KEY_ENTRY_24_5                                                                   (32'h10018a94)
`define KV_REG_KEY_ENTRY_24_5                                                                       (32'ha94)
`define CLP_KV_REG_KEY_ENTRY_24_6                                                                   (32'h10018a98)
`define KV_REG_KEY_ENTRY_24_6                                                                       (32'ha98)
`define CLP_KV_REG_KEY_ENTRY_24_7                                                                   (32'h10018a9c)
`define KV_REG_KEY_ENTRY_24_7                                                                       (32'ha9c)
`define CLP_KV_REG_KEY_ENTRY_24_8                                                                   (32'h10018aa0)
`define KV_REG_KEY_ENTRY_24_8                                                                       (32'haa0)
`define CLP_KV_REG_KEY_ENTRY_24_9                                                                   (32'h10018aa4)
`define KV_REG_KEY_ENTRY_24_9                                                                       (32'haa4)
`define CLP_KV_REG_KEY_ENTRY_24_10                                                                  (32'h10018aa8)
`define KV_REG_KEY_ENTRY_24_10                                                                      (32'haa8)
`define CLP_KV_REG_KEY_ENTRY_24_11                                                                  (32'h10018aac)
`define KV_REG_KEY_ENTRY_24_11                                                                      (32'haac)
`define CLP_KV_REG_KEY_ENTRY_25_0                                                                   (32'h10018ab0)
`define KV_REG_KEY_ENTRY_25_0                                                                       (32'hab0)
`define CLP_KV_REG_KEY_ENTRY_25_1                                                                   (32'h10018ab4)
`define KV_REG_KEY_ENTRY_25_1                                                                       (32'hab4)
`define CLP_KV_REG_KEY_ENTRY_25_2                                                                   (32'h10018ab8)
`define KV_REG_KEY_ENTRY_25_2                                                                       (32'hab8)
`define CLP_KV_REG_KEY_ENTRY_25_3                                                                   (32'h10018abc)
`define KV_REG_KEY_ENTRY_25_3                                                                       (32'habc)
`define CLP_KV_REG_KEY_ENTRY_25_4                                                                   (32'h10018ac0)
`define KV_REG_KEY_ENTRY_25_4                                                                       (32'hac0)
`define CLP_KV_REG_KEY_ENTRY_25_5                                                                   (32'h10018ac4)
`define KV_REG_KEY_ENTRY_25_5                                                                       (32'hac4)
`define CLP_KV_REG_KEY_ENTRY_25_6                                                                   (32'h10018ac8)
`define KV_REG_KEY_ENTRY_25_6                                                                       (32'hac8)
`define CLP_KV_REG_KEY_ENTRY_25_7                                                                   (32'h10018acc)
`define KV_REG_KEY_ENTRY_25_7                                                                       (32'hacc)
`define CLP_KV_REG_KEY_ENTRY_25_8                                                                   (32'h10018ad0)
`define KV_REG_KEY_ENTRY_25_8                                                                       (32'had0)
`define CLP_KV_REG_KEY_ENTRY_25_9                                                                   (32'h10018ad4)
`define KV_REG_KEY_ENTRY_25_9                                                                       (32'had4)
`define CLP_KV_REG_KEY_ENTRY_25_10                                                                  (32'h10018ad8)
`define KV_REG_KEY_ENTRY_25_10                                                                      (32'had8)
`define CLP_KV_REG_KEY_ENTRY_25_11                                                                  (32'h10018adc)
`define KV_REG_KEY_ENTRY_25_11                                                                      (32'hadc)
`define CLP_KV_REG_KEY_ENTRY_26_0                                                                   (32'h10018ae0)
`define KV_REG_KEY_ENTRY_26_0                                                                       (32'hae0)
`define CLP_KV_REG_KEY_ENTRY_26_1                                                                   (32'h10018ae4)
`define KV_REG_KEY_ENTRY_26_1                                                                       (32'hae4)
`define CLP_KV_REG_KEY_ENTRY_26_2                                                                   (32'h10018ae8)
`define KV_REG_KEY_ENTRY_26_2                                                                       (32'hae8)
`define CLP_KV_REG_KEY_ENTRY_26_3                                                                   (32'h10018aec)
`define KV_REG_KEY_ENTRY_26_3                                                                       (32'haec)
`define CLP_KV_REG_KEY_ENTRY_26_4                                                                   (32'h10018af0)
`define KV_REG_KEY_ENTRY_26_4                                                                       (32'haf0)
`define CLP_KV_REG_KEY_ENTRY_26_5                                                                   (32'h10018af4)
`define KV_REG_KEY_ENTRY_26_5                                                                       (32'haf4)
`define CLP_KV_REG_KEY_ENTRY_26_6                                                                   (32'h10018af8)
`define KV_REG_KEY_ENTRY_26_6                                                                       (32'haf8)
`define CLP_KV_REG_KEY_ENTRY_26_7                                                                   (32'h10018afc)
`define KV_REG_KEY_ENTRY_26_7                                                                       (32'hafc)
`define CLP_KV_REG_KEY_ENTRY_26_8                                                                   (32'h10018b00)
`define KV_REG_KEY_ENTRY_26_8                                                                       (32'hb00)
`define CLP_KV_REG_KEY_ENTRY_26_9                                                                   (32'h10018b04)
`define KV_REG_KEY_ENTRY_26_9                                                                       (32'hb04)
`define CLP_KV_REG_KEY_ENTRY_26_10                                                                  (32'h10018b08)
`define KV_REG_KEY_ENTRY_26_10                                                                      (32'hb08)
`define CLP_KV_REG_KEY_ENTRY_26_11                                                                  (32'h10018b0c)
`define KV_REG_KEY_ENTRY_26_11                                                                      (32'hb0c)
`define CLP_KV_REG_KEY_ENTRY_27_0                                                                   (32'h10018b10)
`define KV_REG_KEY_ENTRY_27_0                                                                       (32'hb10)
`define CLP_KV_REG_KEY_ENTRY_27_1                                                                   (32'h10018b14)
`define KV_REG_KEY_ENTRY_27_1                                                                       (32'hb14)
`define CLP_KV_REG_KEY_ENTRY_27_2                                                                   (32'h10018b18)
`define KV_REG_KEY_ENTRY_27_2                                                                       (32'hb18)
`define CLP_KV_REG_KEY_ENTRY_27_3                                                                   (32'h10018b1c)
`define KV_REG_KEY_ENTRY_27_3                                                                       (32'hb1c)
`define CLP_KV_REG_KEY_ENTRY_27_4                                                                   (32'h10018b20)
`define KV_REG_KEY_ENTRY_27_4                                                                       (32'hb20)
`define CLP_KV_REG_KEY_ENTRY_27_5                                                                   (32'h10018b24)
`define KV_REG_KEY_ENTRY_27_5                                                                       (32'hb24)
`define CLP_KV_REG_KEY_ENTRY_27_6                                                                   (32'h10018b28)
`define KV_REG_KEY_ENTRY_27_6                                                                       (32'hb28)
`define CLP_KV_REG_KEY_ENTRY_27_7                                                                   (32'h10018b2c)
`define KV_REG_KEY_ENTRY_27_7                                                                       (32'hb2c)
`define CLP_KV_REG_KEY_ENTRY_27_8                                                                   (32'h10018b30)
`define KV_REG_KEY_ENTRY_27_8                                                                       (32'hb30)
`define CLP_KV_REG_KEY_ENTRY_27_9                                                                   (32'h10018b34)
`define KV_REG_KEY_ENTRY_27_9                                                                       (32'hb34)
`define CLP_KV_REG_KEY_ENTRY_27_10                                                                  (32'h10018b38)
`define KV_REG_KEY_ENTRY_27_10                                                                      (32'hb38)
`define CLP_KV_REG_KEY_ENTRY_27_11                                                                  (32'h10018b3c)
`define KV_REG_KEY_ENTRY_27_11                                                                      (32'hb3c)
`define CLP_KV_REG_KEY_ENTRY_28_0                                                                   (32'h10018b40)
`define KV_REG_KEY_ENTRY_28_0                                                                       (32'hb40)
`define CLP_KV_REG_KEY_ENTRY_28_1                                                                   (32'h10018b44)
`define KV_REG_KEY_ENTRY_28_1                                                                       (32'hb44)
`define CLP_KV_REG_KEY_ENTRY_28_2                                                                   (32'h10018b48)
`define KV_REG_KEY_ENTRY_28_2                                                                       (32'hb48)
`define CLP_KV_REG_KEY_ENTRY_28_3                                                                   (32'h10018b4c)
`define KV_REG_KEY_ENTRY_28_3                                                                       (32'hb4c)
`define CLP_KV_REG_KEY_ENTRY_28_4                                                                   (32'h10018b50)
`define KV_REG_KEY_ENTRY_28_4                                                                       (32'hb50)
`define CLP_KV_REG_KEY_ENTRY_28_5                                                                   (32'h10018b54)
`define KV_REG_KEY_ENTRY_28_5                                                                       (32'hb54)
`define CLP_KV_REG_KEY_ENTRY_28_6                                                                   (32'h10018b58)
`define KV_REG_KEY_ENTRY_28_6                                                                       (32'hb58)
`define CLP_KV_REG_KEY_ENTRY_28_7                                                                   (32'h10018b5c)
`define KV_REG_KEY_ENTRY_28_7                                                                       (32'hb5c)
`define CLP_KV_REG_KEY_ENTRY_28_8                                                                   (32'h10018b60)
`define KV_REG_KEY_ENTRY_28_8                                                                       (32'hb60)
`define CLP_KV_REG_KEY_ENTRY_28_9                                                                   (32'h10018b64)
`define KV_REG_KEY_ENTRY_28_9                                                                       (32'hb64)
`define CLP_KV_REG_KEY_ENTRY_28_10                                                                  (32'h10018b68)
`define KV_REG_KEY_ENTRY_28_10                                                                      (32'hb68)
`define CLP_KV_REG_KEY_ENTRY_28_11                                                                  (32'h10018b6c)
`define KV_REG_KEY_ENTRY_28_11                                                                      (32'hb6c)
`define CLP_KV_REG_KEY_ENTRY_29_0                                                                   (32'h10018b70)
`define KV_REG_KEY_ENTRY_29_0                                                                       (32'hb70)
`define CLP_KV_REG_KEY_ENTRY_29_1                                                                   (32'h10018b74)
`define KV_REG_KEY_ENTRY_29_1                                                                       (32'hb74)
`define CLP_KV_REG_KEY_ENTRY_29_2                                                                   (32'h10018b78)
`define KV_REG_KEY_ENTRY_29_2                                                                       (32'hb78)
`define CLP_KV_REG_KEY_ENTRY_29_3                                                                   (32'h10018b7c)
`define KV_REG_KEY_ENTRY_29_3                                                                       (32'hb7c)
`define CLP_KV_REG_KEY_ENTRY_29_4                                                                   (32'h10018b80)
`define KV_REG_KEY_ENTRY_29_4                                                                       (32'hb80)
`define CLP_KV_REG_KEY_ENTRY_29_5                                                                   (32'h10018b84)
`define KV_REG_KEY_ENTRY_29_5                                                                       (32'hb84)
`define CLP_KV_REG_KEY_ENTRY_29_6                                                                   (32'h10018b88)
`define KV_REG_KEY_ENTRY_29_6                                                                       (32'hb88)
`define CLP_KV_REG_KEY_ENTRY_29_7                                                                   (32'h10018b8c)
`define KV_REG_KEY_ENTRY_29_7                                                                       (32'hb8c)
`define CLP_KV_REG_KEY_ENTRY_29_8                                                                   (32'h10018b90)
`define KV_REG_KEY_ENTRY_29_8                                                                       (32'hb90)
`define CLP_KV_REG_KEY_ENTRY_29_9                                                                   (32'h10018b94)
`define KV_REG_KEY_ENTRY_29_9                                                                       (32'hb94)
`define CLP_KV_REG_KEY_ENTRY_29_10                                                                  (32'h10018b98)
`define KV_REG_KEY_ENTRY_29_10                                                                      (32'hb98)
`define CLP_KV_REG_KEY_ENTRY_29_11                                                                  (32'h10018b9c)
`define KV_REG_KEY_ENTRY_29_11                                                                      (32'hb9c)
`define CLP_KV_REG_KEY_ENTRY_30_0                                                                   (32'h10018ba0)
`define KV_REG_KEY_ENTRY_30_0                                                                       (32'hba0)
`define CLP_KV_REG_KEY_ENTRY_30_1                                                                   (32'h10018ba4)
`define KV_REG_KEY_ENTRY_30_1                                                                       (32'hba4)
`define CLP_KV_REG_KEY_ENTRY_30_2                                                                   (32'h10018ba8)
`define KV_REG_KEY_ENTRY_30_2                                                                       (32'hba8)
`define CLP_KV_REG_KEY_ENTRY_30_3                                                                   (32'h10018bac)
`define KV_REG_KEY_ENTRY_30_3                                                                       (32'hbac)
`define CLP_KV_REG_KEY_ENTRY_30_4                                                                   (32'h10018bb0)
`define KV_REG_KEY_ENTRY_30_4                                                                       (32'hbb0)
`define CLP_KV_REG_KEY_ENTRY_30_5                                                                   (32'h10018bb4)
`define KV_REG_KEY_ENTRY_30_5                                                                       (32'hbb4)
`define CLP_KV_REG_KEY_ENTRY_30_6                                                                   (32'h10018bb8)
`define KV_REG_KEY_ENTRY_30_6                                                                       (32'hbb8)
`define CLP_KV_REG_KEY_ENTRY_30_7                                                                   (32'h10018bbc)
`define KV_REG_KEY_ENTRY_30_7                                                                       (32'hbbc)
`define CLP_KV_REG_KEY_ENTRY_30_8                                                                   (32'h10018bc0)
`define KV_REG_KEY_ENTRY_30_8                                                                       (32'hbc0)
`define CLP_KV_REG_KEY_ENTRY_30_9                                                                   (32'h10018bc4)
`define KV_REG_KEY_ENTRY_30_9                                                                       (32'hbc4)
`define CLP_KV_REG_KEY_ENTRY_30_10                                                                  (32'h10018bc8)
`define KV_REG_KEY_ENTRY_30_10                                                                      (32'hbc8)
`define CLP_KV_REG_KEY_ENTRY_30_11                                                                  (32'h10018bcc)
`define KV_REG_KEY_ENTRY_30_11                                                                      (32'hbcc)
`define CLP_KV_REG_KEY_ENTRY_31_0                                                                   (32'h10018bd0)
`define KV_REG_KEY_ENTRY_31_0                                                                       (32'hbd0)
`define CLP_KV_REG_KEY_ENTRY_31_1                                                                   (32'h10018bd4)
`define KV_REG_KEY_ENTRY_31_1                                                                       (32'hbd4)
`define CLP_KV_REG_KEY_ENTRY_31_2                                                                   (32'h10018bd8)
`define KV_REG_KEY_ENTRY_31_2                                                                       (32'hbd8)
`define CLP_KV_REG_KEY_ENTRY_31_3                                                                   (32'h10018bdc)
`define KV_REG_KEY_ENTRY_31_3                                                                       (32'hbdc)
`define CLP_KV_REG_KEY_ENTRY_31_4                                                                   (32'h10018be0)
`define KV_REG_KEY_ENTRY_31_4                                                                       (32'hbe0)
`define CLP_KV_REG_KEY_ENTRY_31_5                                                                   (32'h10018be4)
`define KV_REG_KEY_ENTRY_31_5                                                                       (32'hbe4)
`define CLP_KV_REG_KEY_ENTRY_31_6                                                                   (32'h10018be8)
`define KV_REG_KEY_ENTRY_31_6                                                                       (32'hbe8)
`define CLP_KV_REG_KEY_ENTRY_31_7                                                                   (32'h10018bec)
`define KV_REG_KEY_ENTRY_31_7                                                                       (32'hbec)
`define CLP_KV_REG_KEY_ENTRY_31_8                                                                   (32'h10018bf0)
`define KV_REG_KEY_ENTRY_31_8                                                                       (32'hbf0)
`define CLP_KV_REG_KEY_ENTRY_31_9                                                                   (32'h10018bf4)
`define KV_REG_KEY_ENTRY_31_9                                                                       (32'hbf4)
`define CLP_KV_REG_KEY_ENTRY_31_10                                                                  (32'h10018bf8)
`define KV_REG_KEY_ENTRY_31_10                                                                      (32'hbf8)
`define CLP_KV_REG_KEY_ENTRY_31_11                                                                  (32'h10018bfc)
`define KV_REG_KEY_ENTRY_31_11                                                                      (32'hbfc)
`define CLP_KV_REG_CLEAR_SECRETS                                                                    (32'h10018c00)
`define KV_REG_CLEAR_SECRETS                                                                        (32'hc00)
`define KV_REG_CLEAR_SECRETS_WR_DEBUG_VALUES_LOW                                                    (0)
`define KV_REG_CLEAR_SECRETS_WR_DEBUG_VALUES_MASK                                                   (32'h1)
`define KV_REG_CLEAR_SECRETS_SEL_DEBUG_VALUE_LOW                                                    (1)
`define KV_REG_CLEAR_SECRETS_SEL_DEBUG_VALUE_MASK                                                   (32'h2)
`define CLP_PV_REG_BASE_ADDR                                                                        (32'h1001a000)
`define CLP_PV_REG_PCR_CTRL_0                                                                       (32'h1001a000)
`define PV_REG_PCR_CTRL_0                                                                           (32'h0)
`define PV_REG_PCR_CTRL_0_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_0_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_0_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_0_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_0_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_0_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_0_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_0_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_1                                                                       (32'h1001a004)
`define PV_REG_PCR_CTRL_1                                                                           (32'h4)
`define PV_REG_PCR_CTRL_1_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_1_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_1_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_1_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_1_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_1_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_1_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_1_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_2                                                                       (32'h1001a008)
`define PV_REG_PCR_CTRL_2                                                                           (32'h8)
`define PV_REG_PCR_CTRL_2_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_2_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_2_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_2_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_2_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_2_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_2_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_2_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_3                                                                       (32'h1001a00c)
`define PV_REG_PCR_CTRL_3                                                                           (32'hc)
`define PV_REG_PCR_CTRL_3_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_3_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_3_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_3_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_3_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_3_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_3_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_3_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_4                                                                       (32'h1001a010)
`define PV_REG_PCR_CTRL_4                                                                           (32'h10)
`define PV_REG_PCR_CTRL_4_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_4_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_4_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_4_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_4_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_4_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_4_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_4_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_5                                                                       (32'h1001a014)
`define PV_REG_PCR_CTRL_5                                                                           (32'h14)
`define PV_REG_PCR_CTRL_5_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_5_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_5_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_5_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_5_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_5_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_5_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_5_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_6                                                                       (32'h1001a018)
`define PV_REG_PCR_CTRL_6                                                                           (32'h18)
`define PV_REG_PCR_CTRL_6_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_6_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_6_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_6_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_6_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_6_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_6_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_6_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_7                                                                       (32'h1001a01c)
`define PV_REG_PCR_CTRL_7                                                                           (32'h1c)
`define PV_REG_PCR_CTRL_7_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_7_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_7_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_7_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_7_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_7_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_7_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_7_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_8                                                                       (32'h1001a020)
`define PV_REG_PCR_CTRL_8                                                                           (32'h20)
`define PV_REG_PCR_CTRL_8_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_8_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_8_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_8_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_8_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_8_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_8_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_8_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_9                                                                       (32'h1001a024)
`define PV_REG_PCR_CTRL_9                                                                           (32'h24)
`define PV_REG_PCR_CTRL_9_LOCK_LOW                                                                  (0)
`define PV_REG_PCR_CTRL_9_LOCK_MASK                                                                 (32'h1)
`define PV_REG_PCR_CTRL_9_CLEAR_LOW                                                                 (1)
`define PV_REG_PCR_CTRL_9_CLEAR_MASK                                                                (32'h2)
`define PV_REG_PCR_CTRL_9_RSVD0_LOW                                                                 (2)
`define PV_REG_PCR_CTRL_9_RSVD0_MASK                                                                (32'h4)
`define PV_REG_PCR_CTRL_9_RSVD1_LOW                                                                 (3)
`define PV_REG_PCR_CTRL_9_RSVD1_MASK                                                                (32'hf8)
`define CLP_PV_REG_PCR_CTRL_10                                                                      (32'h1001a028)
`define PV_REG_PCR_CTRL_10                                                                          (32'h28)
`define PV_REG_PCR_CTRL_10_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_10_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_10_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_10_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_10_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_10_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_10_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_10_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_11                                                                      (32'h1001a02c)
`define PV_REG_PCR_CTRL_11                                                                          (32'h2c)
`define PV_REG_PCR_CTRL_11_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_11_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_11_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_11_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_11_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_11_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_11_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_11_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_12                                                                      (32'h1001a030)
`define PV_REG_PCR_CTRL_12                                                                          (32'h30)
`define PV_REG_PCR_CTRL_12_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_12_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_12_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_12_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_12_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_12_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_12_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_12_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_13                                                                      (32'h1001a034)
`define PV_REG_PCR_CTRL_13                                                                          (32'h34)
`define PV_REG_PCR_CTRL_13_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_13_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_13_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_13_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_13_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_13_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_13_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_13_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_14                                                                      (32'h1001a038)
`define PV_REG_PCR_CTRL_14                                                                          (32'h38)
`define PV_REG_PCR_CTRL_14_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_14_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_14_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_14_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_14_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_14_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_14_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_14_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_15                                                                      (32'h1001a03c)
`define PV_REG_PCR_CTRL_15                                                                          (32'h3c)
`define PV_REG_PCR_CTRL_15_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_15_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_15_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_15_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_15_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_15_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_15_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_15_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_16                                                                      (32'h1001a040)
`define PV_REG_PCR_CTRL_16                                                                          (32'h40)
`define PV_REG_PCR_CTRL_16_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_16_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_16_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_16_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_16_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_16_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_16_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_16_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_17                                                                      (32'h1001a044)
`define PV_REG_PCR_CTRL_17                                                                          (32'h44)
`define PV_REG_PCR_CTRL_17_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_17_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_17_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_17_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_17_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_17_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_17_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_17_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_18                                                                      (32'h1001a048)
`define PV_REG_PCR_CTRL_18                                                                          (32'h48)
`define PV_REG_PCR_CTRL_18_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_18_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_18_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_18_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_18_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_18_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_18_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_18_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_19                                                                      (32'h1001a04c)
`define PV_REG_PCR_CTRL_19                                                                          (32'h4c)
`define PV_REG_PCR_CTRL_19_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_19_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_19_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_19_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_19_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_19_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_19_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_19_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_20                                                                      (32'h1001a050)
`define PV_REG_PCR_CTRL_20                                                                          (32'h50)
`define PV_REG_PCR_CTRL_20_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_20_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_20_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_20_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_20_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_20_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_20_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_20_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_21                                                                      (32'h1001a054)
`define PV_REG_PCR_CTRL_21                                                                          (32'h54)
`define PV_REG_PCR_CTRL_21_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_21_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_21_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_21_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_21_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_21_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_21_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_21_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_22                                                                      (32'h1001a058)
`define PV_REG_PCR_CTRL_22                                                                          (32'h58)
`define PV_REG_PCR_CTRL_22_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_22_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_22_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_22_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_22_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_22_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_22_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_22_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_23                                                                      (32'h1001a05c)
`define PV_REG_PCR_CTRL_23                                                                          (32'h5c)
`define PV_REG_PCR_CTRL_23_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_23_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_23_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_23_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_23_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_23_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_23_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_23_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_24                                                                      (32'h1001a060)
`define PV_REG_PCR_CTRL_24                                                                          (32'h60)
`define PV_REG_PCR_CTRL_24_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_24_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_24_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_24_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_24_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_24_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_24_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_24_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_25                                                                      (32'h1001a064)
`define PV_REG_PCR_CTRL_25                                                                          (32'h64)
`define PV_REG_PCR_CTRL_25_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_25_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_25_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_25_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_25_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_25_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_25_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_25_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_26                                                                      (32'h1001a068)
`define PV_REG_PCR_CTRL_26                                                                          (32'h68)
`define PV_REG_PCR_CTRL_26_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_26_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_26_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_26_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_26_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_26_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_26_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_26_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_27                                                                      (32'h1001a06c)
`define PV_REG_PCR_CTRL_27                                                                          (32'h6c)
`define PV_REG_PCR_CTRL_27_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_27_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_27_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_27_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_27_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_27_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_27_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_27_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_28                                                                      (32'h1001a070)
`define PV_REG_PCR_CTRL_28                                                                          (32'h70)
`define PV_REG_PCR_CTRL_28_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_28_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_28_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_28_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_28_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_28_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_28_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_28_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_29                                                                      (32'h1001a074)
`define PV_REG_PCR_CTRL_29                                                                          (32'h74)
`define PV_REG_PCR_CTRL_29_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_29_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_29_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_29_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_29_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_29_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_29_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_29_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_30                                                                      (32'h1001a078)
`define PV_REG_PCR_CTRL_30                                                                          (32'h78)
`define PV_REG_PCR_CTRL_30_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_30_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_30_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_30_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_30_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_30_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_30_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_30_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_CTRL_31                                                                      (32'h1001a07c)
`define PV_REG_PCR_CTRL_31                                                                          (32'h7c)
`define PV_REG_PCR_CTRL_31_LOCK_LOW                                                                 (0)
`define PV_REG_PCR_CTRL_31_LOCK_MASK                                                                (32'h1)
`define PV_REG_PCR_CTRL_31_CLEAR_LOW                                                                (1)
`define PV_REG_PCR_CTRL_31_CLEAR_MASK                                                               (32'h2)
`define PV_REG_PCR_CTRL_31_RSVD0_LOW                                                                (2)
`define PV_REG_PCR_CTRL_31_RSVD0_MASK                                                               (32'h4)
`define PV_REG_PCR_CTRL_31_RSVD1_LOW                                                                (3)
`define PV_REG_PCR_CTRL_31_RSVD1_MASK                                                               (32'hf8)
`define CLP_PV_REG_PCR_ENTRY_0_0                                                                    (32'h1001a600)
`define PV_REG_PCR_ENTRY_0_0                                                                        (32'h600)
`define CLP_PV_REG_PCR_ENTRY_0_1                                                                    (32'h1001a604)
`define PV_REG_PCR_ENTRY_0_1                                                                        (32'h604)
`define CLP_PV_REG_PCR_ENTRY_0_2                                                                    (32'h1001a608)
`define PV_REG_PCR_ENTRY_0_2                                                                        (32'h608)
`define CLP_PV_REG_PCR_ENTRY_0_3                                                                    (32'h1001a60c)
`define PV_REG_PCR_ENTRY_0_3                                                                        (32'h60c)
`define CLP_PV_REG_PCR_ENTRY_0_4                                                                    (32'h1001a610)
`define PV_REG_PCR_ENTRY_0_4                                                                        (32'h610)
`define CLP_PV_REG_PCR_ENTRY_0_5                                                                    (32'h1001a614)
`define PV_REG_PCR_ENTRY_0_5                                                                        (32'h614)
`define CLP_PV_REG_PCR_ENTRY_0_6                                                                    (32'h1001a618)
`define PV_REG_PCR_ENTRY_0_6                                                                        (32'h618)
`define CLP_PV_REG_PCR_ENTRY_0_7                                                                    (32'h1001a61c)
`define PV_REG_PCR_ENTRY_0_7                                                                        (32'h61c)
`define CLP_PV_REG_PCR_ENTRY_0_8                                                                    (32'h1001a620)
`define PV_REG_PCR_ENTRY_0_8                                                                        (32'h620)
`define CLP_PV_REG_PCR_ENTRY_0_9                                                                    (32'h1001a624)
`define PV_REG_PCR_ENTRY_0_9                                                                        (32'h624)
`define CLP_PV_REG_PCR_ENTRY_0_10                                                                   (32'h1001a628)
`define PV_REG_PCR_ENTRY_0_10                                                                       (32'h628)
`define CLP_PV_REG_PCR_ENTRY_0_11                                                                   (32'h1001a62c)
`define PV_REG_PCR_ENTRY_0_11                                                                       (32'h62c)
`define CLP_PV_REG_PCR_ENTRY_1_0                                                                    (32'h1001a630)
`define PV_REG_PCR_ENTRY_1_0                                                                        (32'h630)
`define CLP_PV_REG_PCR_ENTRY_1_1                                                                    (32'h1001a634)
`define PV_REG_PCR_ENTRY_1_1                                                                        (32'h634)
`define CLP_PV_REG_PCR_ENTRY_1_2                                                                    (32'h1001a638)
`define PV_REG_PCR_ENTRY_1_2                                                                        (32'h638)
`define CLP_PV_REG_PCR_ENTRY_1_3                                                                    (32'h1001a63c)
`define PV_REG_PCR_ENTRY_1_3                                                                        (32'h63c)
`define CLP_PV_REG_PCR_ENTRY_1_4                                                                    (32'h1001a640)
`define PV_REG_PCR_ENTRY_1_4                                                                        (32'h640)
`define CLP_PV_REG_PCR_ENTRY_1_5                                                                    (32'h1001a644)
`define PV_REG_PCR_ENTRY_1_5                                                                        (32'h644)
`define CLP_PV_REG_PCR_ENTRY_1_6                                                                    (32'h1001a648)
`define PV_REG_PCR_ENTRY_1_6                                                                        (32'h648)
`define CLP_PV_REG_PCR_ENTRY_1_7                                                                    (32'h1001a64c)
`define PV_REG_PCR_ENTRY_1_7                                                                        (32'h64c)
`define CLP_PV_REG_PCR_ENTRY_1_8                                                                    (32'h1001a650)
`define PV_REG_PCR_ENTRY_1_8                                                                        (32'h650)
`define CLP_PV_REG_PCR_ENTRY_1_9                                                                    (32'h1001a654)
`define PV_REG_PCR_ENTRY_1_9                                                                        (32'h654)
`define CLP_PV_REG_PCR_ENTRY_1_10                                                                   (32'h1001a658)
`define PV_REG_PCR_ENTRY_1_10                                                                       (32'h658)
`define CLP_PV_REG_PCR_ENTRY_1_11                                                                   (32'h1001a65c)
`define PV_REG_PCR_ENTRY_1_11                                                                       (32'h65c)
`define CLP_PV_REG_PCR_ENTRY_2_0                                                                    (32'h1001a660)
`define PV_REG_PCR_ENTRY_2_0                                                                        (32'h660)
`define CLP_PV_REG_PCR_ENTRY_2_1                                                                    (32'h1001a664)
`define PV_REG_PCR_ENTRY_2_1                                                                        (32'h664)
`define CLP_PV_REG_PCR_ENTRY_2_2                                                                    (32'h1001a668)
`define PV_REG_PCR_ENTRY_2_2                                                                        (32'h668)
`define CLP_PV_REG_PCR_ENTRY_2_3                                                                    (32'h1001a66c)
`define PV_REG_PCR_ENTRY_2_3                                                                        (32'h66c)
`define CLP_PV_REG_PCR_ENTRY_2_4                                                                    (32'h1001a670)
`define PV_REG_PCR_ENTRY_2_4                                                                        (32'h670)
`define CLP_PV_REG_PCR_ENTRY_2_5                                                                    (32'h1001a674)
`define PV_REG_PCR_ENTRY_2_5                                                                        (32'h674)
`define CLP_PV_REG_PCR_ENTRY_2_6                                                                    (32'h1001a678)
`define PV_REG_PCR_ENTRY_2_6                                                                        (32'h678)
`define CLP_PV_REG_PCR_ENTRY_2_7                                                                    (32'h1001a67c)
`define PV_REG_PCR_ENTRY_2_7                                                                        (32'h67c)
`define CLP_PV_REG_PCR_ENTRY_2_8                                                                    (32'h1001a680)
`define PV_REG_PCR_ENTRY_2_8                                                                        (32'h680)
`define CLP_PV_REG_PCR_ENTRY_2_9                                                                    (32'h1001a684)
`define PV_REG_PCR_ENTRY_2_9                                                                        (32'h684)
`define CLP_PV_REG_PCR_ENTRY_2_10                                                                   (32'h1001a688)
`define PV_REG_PCR_ENTRY_2_10                                                                       (32'h688)
`define CLP_PV_REG_PCR_ENTRY_2_11                                                                   (32'h1001a68c)
`define PV_REG_PCR_ENTRY_2_11                                                                       (32'h68c)
`define CLP_PV_REG_PCR_ENTRY_3_0                                                                    (32'h1001a690)
`define PV_REG_PCR_ENTRY_3_0                                                                        (32'h690)
`define CLP_PV_REG_PCR_ENTRY_3_1                                                                    (32'h1001a694)
`define PV_REG_PCR_ENTRY_3_1                                                                        (32'h694)
`define CLP_PV_REG_PCR_ENTRY_3_2                                                                    (32'h1001a698)
`define PV_REG_PCR_ENTRY_3_2                                                                        (32'h698)
`define CLP_PV_REG_PCR_ENTRY_3_3                                                                    (32'h1001a69c)
`define PV_REG_PCR_ENTRY_3_3                                                                        (32'h69c)
`define CLP_PV_REG_PCR_ENTRY_3_4                                                                    (32'h1001a6a0)
`define PV_REG_PCR_ENTRY_3_4                                                                        (32'h6a0)
`define CLP_PV_REG_PCR_ENTRY_3_5                                                                    (32'h1001a6a4)
`define PV_REG_PCR_ENTRY_3_5                                                                        (32'h6a4)
`define CLP_PV_REG_PCR_ENTRY_3_6                                                                    (32'h1001a6a8)
`define PV_REG_PCR_ENTRY_3_6                                                                        (32'h6a8)
`define CLP_PV_REG_PCR_ENTRY_3_7                                                                    (32'h1001a6ac)
`define PV_REG_PCR_ENTRY_3_7                                                                        (32'h6ac)
`define CLP_PV_REG_PCR_ENTRY_3_8                                                                    (32'h1001a6b0)
`define PV_REG_PCR_ENTRY_3_8                                                                        (32'h6b0)
`define CLP_PV_REG_PCR_ENTRY_3_9                                                                    (32'h1001a6b4)
`define PV_REG_PCR_ENTRY_3_9                                                                        (32'h6b4)
`define CLP_PV_REG_PCR_ENTRY_3_10                                                                   (32'h1001a6b8)
`define PV_REG_PCR_ENTRY_3_10                                                                       (32'h6b8)
`define CLP_PV_REG_PCR_ENTRY_3_11                                                                   (32'h1001a6bc)
`define PV_REG_PCR_ENTRY_3_11                                                                       (32'h6bc)
`define CLP_PV_REG_PCR_ENTRY_4_0                                                                    (32'h1001a6c0)
`define PV_REG_PCR_ENTRY_4_0                                                                        (32'h6c0)
`define CLP_PV_REG_PCR_ENTRY_4_1                                                                    (32'h1001a6c4)
`define PV_REG_PCR_ENTRY_4_1                                                                        (32'h6c4)
`define CLP_PV_REG_PCR_ENTRY_4_2                                                                    (32'h1001a6c8)
`define PV_REG_PCR_ENTRY_4_2                                                                        (32'h6c8)
`define CLP_PV_REG_PCR_ENTRY_4_3                                                                    (32'h1001a6cc)
`define PV_REG_PCR_ENTRY_4_3                                                                        (32'h6cc)
`define CLP_PV_REG_PCR_ENTRY_4_4                                                                    (32'h1001a6d0)
`define PV_REG_PCR_ENTRY_4_4                                                                        (32'h6d0)
`define CLP_PV_REG_PCR_ENTRY_4_5                                                                    (32'h1001a6d4)
`define PV_REG_PCR_ENTRY_4_5                                                                        (32'h6d4)
`define CLP_PV_REG_PCR_ENTRY_4_6                                                                    (32'h1001a6d8)
`define PV_REG_PCR_ENTRY_4_6                                                                        (32'h6d8)
`define CLP_PV_REG_PCR_ENTRY_4_7                                                                    (32'h1001a6dc)
`define PV_REG_PCR_ENTRY_4_7                                                                        (32'h6dc)
`define CLP_PV_REG_PCR_ENTRY_4_8                                                                    (32'h1001a6e0)
`define PV_REG_PCR_ENTRY_4_8                                                                        (32'h6e0)
`define CLP_PV_REG_PCR_ENTRY_4_9                                                                    (32'h1001a6e4)
`define PV_REG_PCR_ENTRY_4_9                                                                        (32'h6e4)
`define CLP_PV_REG_PCR_ENTRY_4_10                                                                   (32'h1001a6e8)
`define PV_REG_PCR_ENTRY_4_10                                                                       (32'h6e8)
`define CLP_PV_REG_PCR_ENTRY_4_11                                                                   (32'h1001a6ec)
`define PV_REG_PCR_ENTRY_4_11                                                                       (32'h6ec)
`define CLP_PV_REG_PCR_ENTRY_5_0                                                                    (32'h1001a6f0)
`define PV_REG_PCR_ENTRY_5_0                                                                        (32'h6f0)
`define CLP_PV_REG_PCR_ENTRY_5_1                                                                    (32'h1001a6f4)
`define PV_REG_PCR_ENTRY_5_1                                                                        (32'h6f4)
`define CLP_PV_REG_PCR_ENTRY_5_2                                                                    (32'h1001a6f8)
`define PV_REG_PCR_ENTRY_5_2                                                                        (32'h6f8)
`define CLP_PV_REG_PCR_ENTRY_5_3                                                                    (32'h1001a6fc)
`define PV_REG_PCR_ENTRY_5_3                                                                        (32'h6fc)
`define CLP_PV_REG_PCR_ENTRY_5_4                                                                    (32'h1001a700)
`define PV_REG_PCR_ENTRY_5_4                                                                        (32'h700)
`define CLP_PV_REG_PCR_ENTRY_5_5                                                                    (32'h1001a704)
`define PV_REG_PCR_ENTRY_5_5                                                                        (32'h704)
`define CLP_PV_REG_PCR_ENTRY_5_6                                                                    (32'h1001a708)
`define PV_REG_PCR_ENTRY_5_6                                                                        (32'h708)
`define CLP_PV_REG_PCR_ENTRY_5_7                                                                    (32'h1001a70c)
`define PV_REG_PCR_ENTRY_5_7                                                                        (32'h70c)
`define CLP_PV_REG_PCR_ENTRY_5_8                                                                    (32'h1001a710)
`define PV_REG_PCR_ENTRY_5_8                                                                        (32'h710)
`define CLP_PV_REG_PCR_ENTRY_5_9                                                                    (32'h1001a714)
`define PV_REG_PCR_ENTRY_5_9                                                                        (32'h714)
`define CLP_PV_REG_PCR_ENTRY_5_10                                                                   (32'h1001a718)
`define PV_REG_PCR_ENTRY_5_10                                                                       (32'h718)
`define CLP_PV_REG_PCR_ENTRY_5_11                                                                   (32'h1001a71c)
`define PV_REG_PCR_ENTRY_5_11                                                                       (32'h71c)
`define CLP_PV_REG_PCR_ENTRY_6_0                                                                    (32'h1001a720)
`define PV_REG_PCR_ENTRY_6_0                                                                        (32'h720)
`define CLP_PV_REG_PCR_ENTRY_6_1                                                                    (32'h1001a724)
`define PV_REG_PCR_ENTRY_6_1                                                                        (32'h724)
`define CLP_PV_REG_PCR_ENTRY_6_2                                                                    (32'h1001a728)
`define PV_REG_PCR_ENTRY_6_2                                                                        (32'h728)
`define CLP_PV_REG_PCR_ENTRY_6_3                                                                    (32'h1001a72c)
`define PV_REG_PCR_ENTRY_6_3                                                                        (32'h72c)
`define CLP_PV_REG_PCR_ENTRY_6_4                                                                    (32'h1001a730)
`define PV_REG_PCR_ENTRY_6_4                                                                        (32'h730)
`define CLP_PV_REG_PCR_ENTRY_6_5                                                                    (32'h1001a734)
`define PV_REG_PCR_ENTRY_6_5                                                                        (32'h734)
`define CLP_PV_REG_PCR_ENTRY_6_6                                                                    (32'h1001a738)
`define PV_REG_PCR_ENTRY_6_6                                                                        (32'h738)
`define CLP_PV_REG_PCR_ENTRY_6_7                                                                    (32'h1001a73c)
`define PV_REG_PCR_ENTRY_6_7                                                                        (32'h73c)
`define CLP_PV_REG_PCR_ENTRY_6_8                                                                    (32'h1001a740)
`define PV_REG_PCR_ENTRY_6_8                                                                        (32'h740)
`define CLP_PV_REG_PCR_ENTRY_6_9                                                                    (32'h1001a744)
`define PV_REG_PCR_ENTRY_6_9                                                                        (32'h744)
`define CLP_PV_REG_PCR_ENTRY_6_10                                                                   (32'h1001a748)
`define PV_REG_PCR_ENTRY_6_10                                                                       (32'h748)
`define CLP_PV_REG_PCR_ENTRY_6_11                                                                   (32'h1001a74c)
`define PV_REG_PCR_ENTRY_6_11                                                                       (32'h74c)
`define CLP_PV_REG_PCR_ENTRY_7_0                                                                    (32'h1001a750)
`define PV_REG_PCR_ENTRY_7_0                                                                        (32'h750)
`define CLP_PV_REG_PCR_ENTRY_7_1                                                                    (32'h1001a754)
`define PV_REG_PCR_ENTRY_7_1                                                                        (32'h754)
`define CLP_PV_REG_PCR_ENTRY_7_2                                                                    (32'h1001a758)
`define PV_REG_PCR_ENTRY_7_2                                                                        (32'h758)
`define CLP_PV_REG_PCR_ENTRY_7_3                                                                    (32'h1001a75c)
`define PV_REG_PCR_ENTRY_7_3                                                                        (32'h75c)
`define CLP_PV_REG_PCR_ENTRY_7_4                                                                    (32'h1001a760)
`define PV_REG_PCR_ENTRY_7_4                                                                        (32'h760)
`define CLP_PV_REG_PCR_ENTRY_7_5                                                                    (32'h1001a764)
`define PV_REG_PCR_ENTRY_7_5                                                                        (32'h764)
`define CLP_PV_REG_PCR_ENTRY_7_6                                                                    (32'h1001a768)
`define PV_REG_PCR_ENTRY_7_6                                                                        (32'h768)
`define CLP_PV_REG_PCR_ENTRY_7_7                                                                    (32'h1001a76c)
`define PV_REG_PCR_ENTRY_7_7                                                                        (32'h76c)
`define CLP_PV_REG_PCR_ENTRY_7_8                                                                    (32'h1001a770)
`define PV_REG_PCR_ENTRY_7_8                                                                        (32'h770)
`define CLP_PV_REG_PCR_ENTRY_7_9                                                                    (32'h1001a774)
`define PV_REG_PCR_ENTRY_7_9                                                                        (32'h774)
`define CLP_PV_REG_PCR_ENTRY_7_10                                                                   (32'h1001a778)
`define PV_REG_PCR_ENTRY_7_10                                                                       (32'h778)
`define CLP_PV_REG_PCR_ENTRY_7_11                                                                   (32'h1001a77c)
`define PV_REG_PCR_ENTRY_7_11                                                                       (32'h77c)
`define CLP_PV_REG_PCR_ENTRY_8_0                                                                    (32'h1001a780)
`define PV_REG_PCR_ENTRY_8_0                                                                        (32'h780)
`define CLP_PV_REG_PCR_ENTRY_8_1                                                                    (32'h1001a784)
`define PV_REG_PCR_ENTRY_8_1                                                                        (32'h784)
`define CLP_PV_REG_PCR_ENTRY_8_2                                                                    (32'h1001a788)
`define PV_REG_PCR_ENTRY_8_2                                                                        (32'h788)
`define CLP_PV_REG_PCR_ENTRY_8_3                                                                    (32'h1001a78c)
`define PV_REG_PCR_ENTRY_8_3                                                                        (32'h78c)
`define CLP_PV_REG_PCR_ENTRY_8_4                                                                    (32'h1001a790)
`define PV_REG_PCR_ENTRY_8_4                                                                        (32'h790)
`define CLP_PV_REG_PCR_ENTRY_8_5                                                                    (32'h1001a794)
`define PV_REG_PCR_ENTRY_8_5                                                                        (32'h794)
`define CLP_PV_REG_PCR_ENTRY_8_6                                                                    (32'h1001a798)
`define PV_REG_PCR_ENTRY_8_6                                                                        (32'h798)
`define CLP_PV_REG_PCR_ENTRY_8_7                                                                    (32'h1001a79c)
`define PV_REG_PCR_ENTRY_8_7                                                                        (32'h79c)
`define CLP_PV_REG_PCR_ENTRY_8_8                                                                    (32'h1001a7a0)
`define PV_REG_PCR_ENTRY_8_8                                                                        (32'h7a0)
`define CLP_PV_REG_PCR_ENTRY_8_9                                                                    (32'h1001a7a4)
`define PV_REG_PCR_ENTRY_8_9                                                                        (32'h7a4)
`define CLP_PV_REG_PCR_ENTRY_8_10                                                                   (32'h1001a7a8)
`define PV_REG_PCR_ENTRY_8_10                                                                       (32'h7a8)
`define CLP_PV_REG_PCR_ENTRY_8_11                                                                   (32'h1001a7ac)
`define PV_REG_PCR_ENTRY_8_11                                                                       (32'h7ac)
`define CLP_PV_REG_PCR_ENTRY_9_0                                                                    (32'h1001a7b0)
`define PV_REG_PCR_ENTRY_9_0                                                                        (32'h7b0)
`define CLP_PV_REG_PCR_ENTRY_9_1                                                                    (32'h1001a7b4)
`define PV_REG_PCR_ENTRY_9_1                                                                        (32'h7b4)
`define CLP_PV_REG_PCR_ENTRY_9_2                                                                    (32'h1001a7b8)
`define PV_REG_PCR_ENTRY_9_2                                                                        (32'h7b8)
`define CLP_PV_REG_PCR_ENTRY_9_3                                                                    (32'h1001a7bc)
`define PV_REG_PCR_ENTRY_9_3                                                                        (32'h7bc)
`define CLP_PV_REG_PCR_ENTRY_9_4                                                                    (32'h1001a7c0)
`define PV_REG_PCR_ENTRY_9_4                                                                        (32'h7c0)
`define CLP_PV_REG_PCR_ENTRY_9_5                                                                    (32'h1001a7c4)
`define PV_REG_PCR_ENTRY_9_5                                                                        (32'h7c4)
`define CLP_PV_REG_PCR_ENTRY_9_6                                                                    (32'h1001a7c8)
`define PV_REG_PCR_ENTRY_9_6                                                                        (32'h7c8)
`define CLP_PV_REG_PCR_ENTRY_9_7                                                                    (32'h1001a7cc)
`define PV_REG_PCR_ENTRY_9_7                                                                        (32'h7cc)
`define CLP_PV_REG_PCR_ENTRY_9_8                                                                    (32'h1001a7d0)
`define PV_REG_PCR_ENTRY_9_8                                                                        (32'h7d0)
`define CLP_PV_REG_PCR_ENTRY_9_9                                                                    (32'h1001a7d4)
`define PV_REG_PCR_ENTRY_9_9                                                                        (32'h7d4)
`define CLP_PV_REG_PCR_ENTRY_9_10                                                                   (32'h1001a7d8)
`define PV_REG_PCR_ENTRY_9_10                                                                       (32'h7d8)
`define CLP_PV_REG_PCR_ENTRY_9_11                                                                   (32'h1001a7dc)
`define PV_REG_PCR_ENTRY_9_11                                                                       (32'h7dc)
`define CLP_PV_REG_PCR_ENTRY_10_0                                                                   (32'h1001a7e0)
`define PV_REG_PCR_ENTRY_10_0                                                                       (32'h7e0)
`define CLP_PV_REG_PCR_ENTRY_10_1                                                                   (32'h1001a7e4)
`define PV_REG_PCR_ENTRY_10_1                                                                       (32'h7e4)
`define CLP_PV_REG_PCR_ENTRY_10_2                                                                   (32'h1001a7e8)
`define PV_REG_PCR_ENTRY_10_2                                                                       (32'h7e8)
`define CLP_PV_REG_PCR_ENTRY_10_3                                                                   (32'h1001a7ec)
`define PV_REG_PCR_ENTRY_10_3                                                                       (32'h7ec)
`define CLP_PV_REG_PCR_ENTRY_10_4                                                                   (32'h1001a7f0)
`define PV_REG_PCR_ENTRY_10_4                                                                       (32'h7f0)
`define CLP_PV_REG_PCR_ENTRY_10_5                                                                   (32'h1001a7f4)
`define PV_REG_PCR_ENTRY_10_5                                                                       (32'h7f4)
`define CLP_PV_REG_PCR_ENTRY_10_6                                                                   (32'h1001a7f8)
`define PV_REG_PCR_ENTRY_10_6                                                                       (32'h7f8)
`define CLP_PV_REG_PCR_ENTRY_10_7                                                                   (32'h1001a7fc)
`define PV_REG_PCR_ENTRY_10_7                                                                       (32'h7fc)
`define CLP_PV_REG_PCR_ENTRY_10_8                                                                   (32'h1001a800)
`define PV_REG_PCR_ENTRY_10_8                                                                       (32'h800)
`define CLP_PV_REG_PCR_ENTRY_10_9                                                                   (32'h1001a804)
`define PV_REG_PCR_ENTRY_10_9                                                                       (32'h804)
`define CLP_PV_REG_PCR_ENTRY_10_10                                                                  (32'h1001a808)
`define PV_REG_PCR_ENTRY_10_10                                                                      (32'h808)
`define CLP_PV_REG_PCR_ENTRY_10_11                                                                  (32'h1001a80c)
`define PV_REG_PCR_ENTRY_10_11                                                                      (32'h80c)
`define CLP_PV_REG_PCR_ENTRY_11_0                                                                   (32'h1001a810)
`define PV_REG_PCR_ENTRY_11_0                                                                       (32'h810)
`define CLP_PV_REG_PCR_ENTRY_11_1                                                                   (32'h1001a814)
`define PV_REG_PCR_ENTRY_11_1                                                                       (32'h814)
`define CLP_PV_REG_PCR_ENTRY_11_2                                                                   (32'h1001a818)
`define PV_REG_PCR_ENTRY_11_2                                                                       (32'h818)
`define CLP_PV_REG_PCR_ENTRY_11_3                                                                   (32'h1001a81c)
`define PV_REG_PCR_ENTRY_11_3                                                                       (32'h81c)
`define CLP_PV_REG_PCR_ENTRY_11_4                                                                   (32'h1001a820)
`define PV_REG_PCR_ENTRY_11_4                                                                       (32'h820)
`define CLP_PV_REG_PCR_ENTRY_11_5                                                                   (32'h1001a824)
`define PV_REG_PCR_ENTRY_11_5                                                                       (32'h824)
`define CLP_PV_REG_PCR_ENTRY_11_6                                                                   (32'h1001a828)
`define PV_REG_PCR_ENTRY_11_6                                                                       (32'h828)
`define CLP_PV_REG_PCR_ENTRY_11_7                                                                   (32'h1001a82c)
`define PV_REG_PCR_ENTRY_11_7                                                                       (32'h82c)
`define CLP_PV_REG_PCR_ENTRY_11_8                                                                   (32'h1001a830)
`define PV_REG_PCR_ENTRY_11_8                                                                       (32'h830)
`define CLP_PV_REG_PCR_ENTRY_11_9                                                                   (32'h1001a834)
`define PV_REG_PCR_ENTRY_11_9                                                                       (32'h834)
`define CLP_PV_REG_PCR_ENTRY_11_10                                                                  (32'h1001a838)
`define PV_REG_PCR_ENTRY_11_10                                                                      (32'h838)
`define CLP_PV_REG_PCR_ENTRY_11_11                                                                  (32'h1001a83c)
`define PV_REG_PCR_ENTRY_11_11                                                                      (32'h83c)
`define CLP_PV_REG_PCR_ENTRY_12_0                                                                   (32'h1001a840)
`define PV_REG_PCR_ENTRY_12_0                                                                       (32'h840)
`define CLP_PV_REG_PCR_ENTRY_12_1                                                                   (32'h1001a844)
`define PV_REG_PCR_ENTRY_12_1                                                                       (32'h844)
`define CLP_PV_REG_PCR_ENTRY_12_2                                                                   (32'h1001a848)
`define PV_REG_PCR_ENTRY_12_2                                                                       (32'h848)
`define CLP_PV_REG_PCR_ENTRY_12_3                                                                   (32'h1001a84c)
`define PV_REG_PCR_ENTRY_12_3                                                                       (32'h84c)
`define CLP_PV_REG_PCR_ENTRY_12_4                                                                   (32'h1001a850)
`define PV_REG_PCR_ENTRY_12_4                                                                       (32'h850)
`define CLP_PV_REG_PCR_ENTRY_12_5                                                                   (32'h1001a854)
`define PV_REG_PCR_ENTRY_12_5                                                                       (32'h854)
`define CLP_PV_REG_PCR_ENTRY_12_6                                                                   (32'h1001a858)
`define PV_REG_PCR_ENTRY_12_6                                                                       (32'h858)
`define CLP_PV_REG_PCR_ENTRY_12_7                                                                   (32'h1001a85c)
`define PV_REG_PCR_ENTRY_12_7                                                                       (32'h85c)
`define CLP_PV_REG_PCR_ENTRY_12_8                                                                   (32'h1001a860)
`define PV_REG_PCR_ENTRY_12_8                                                                       (32'h860)
`define CLP_PV_REG_PCR_ENTRY_12_9                                                                   (32'h1001a864)
`define PV_REG_PCR_ENTRY_12_9                                                                       (32'h864)
`define CLP_PV_REG_PCR_ENTRY_12_10                                                                  (32'h1001a868)
`define PV_REG_PCR_ENTRY_12_10                                                                      (32'h868)
`define CLP_PV_REG_PCR_ENTRY_12_11                                                                  (32'h1001a86c)
`define PV_REG_PCR_ENTRY_12_11                                                                      (32'h86c)
`define CLP_PV_REG_PCR_ENTRY_13_0                                                                   (32'h1001a870)
`define PV_REG_PCR_ENTRY_13_0                                                                       (32'h870)
`define CLP_PV_REG_PCR_ENTRY_13_1                                                                   (32'h1001a874)
`define PV_REG_PCR_ENTRY_13_1                                                                       (32'h874)
`define CLP_PV_REG_PCR_ENTRY_13_2                                                                   (32'h1001a878)
`define PV_REG_PCR_ENTRY_13_2                                                                       (32'h878)
`define CLP_PV_REG_PCR_ENTRY_13_3                                                                   (32'h1001a87c)
`define PV_REG_PCR_ENTRY_13_3                                                                       (32'h87c)
`define CLP_PV_REG_PCR_ENTRY_13_4                                                                   (32'h1001a880)
`define PV_REG_PCR_ENTRY_13_4                                                                       (32'h880)
`define CLP_PV_REG_PCR_ENTRY_13_5                                                                   (32'h1001a884)
`define PV_REG_PCR_ENTRY_13_5                                                                       (32'h884)
`define CLP_PV_REG_PCR_ENTRY_13_6                                                                   (32'h1001a888)
`define PV_REG_PCR_ENTRY_13_6                                                                       (32'h888)
`define CLP_PV_REG_PCR_ENTRY_13_7                                                                   (32'h1001a88c)
`define PV_REG_PCR_ENTRY_13_7                                                                       (32'h88c)
`define CLP_PV_REG_PCR_ENTRY_13_8                                                                   (32'h1001a890)
`define PV_REG_PCR_ENTRY_13_8                                                                       (32'h890)
`define CLP_PV_REG_PCR_ENTRY_13_9                                                                   (32'h1001a894)
`define PV_REG_PCR_ENTRY_13_9                                                                       (32'h894)
`define CLP_PV_REG_PCR_ENTRY_13_10                                                                  (32'h1001a898)
`define PV_REG_PCR_ENTRY_13_10                                                                      (32'h898)
`define CLP_PV_REG_PCR_ENTRY_13_11                                                                  (32'h1001a89c)
`define PV_REG_PCR_ENTRY_13_11                                                                      (32'h89c)
`define CLP_PV_REG_PCR_ENTRY_14_0                                                                   (32'h1001a8a0)
`define PV_REG_PCR_ENTRY_14_0                                                                       (32'h8a0)
`define CLP_PV_REG_PCR_ENTRY_14_1                                                                   (32'h1001a8a4)
`define PV_REG_PCR_ENTRY_14_1                                                                       (32'h8a4)
`define CLP_PV_REG_PCR_ENTRY_14_2                                                                   (32'h1001a8a8)
`define PV_REG_PCR_ENTRY_14_2                                                                       (32'h8a8)
`define CLP_PV_REG_PCR_ENTRY_14_3                                                                   (32'h1001a8ac)
`define PV_REG_PCR_ENTRY_14_3                                                                       (32'h8ac)
`define CLP_PV_REG_PCR_ENTRY_14_4                                                                   (32'h1001a8b0)
`define PV_REG_PCR_ENTRY_14_4                                                                       (32'h8b0)
`define CLP_PV_REG_PCR_ENTRY_14_5                                                                   (32'h1001a8b4)
`define PV_REG_PCR_ENTRY_14_5                                                                       (32'h8b4)
`define CLP_PV_REG_PCR_ENTRY_14_6                                                                   (32'h1001a8b8)
`define PV_REG_PCR_ENTRY_14_6                                                                       (32'h8b8)
`define CLP_PV_REG_PCR_ENTRY_14_7                                                                   (32'h1001a8bc)
`define PV_REG_PCR_ENTRY_14_7                                                                       (32'h8bc)
`define CLP_PV_REG_PCR_ENTRY_14_8                                                                   (32'h1001a8c0)
`define PV_REG_PCR_ENTRY_14_8                                                                       (32'h8c0)
`define CLP_PV_REG_PCR_ENTRY_14_9                                                                   (32'h1001a8c4)
`define PV_REG_PCR_ENTRY_14_9                                                                       (32'h8c4)
`define CLP_PV_REG_PCR_ENTRY_14_10                                                                  (32'h1001a8c8)
`define PV_REG_PCR_ENTRY_14_10                                                                      (32'h8c8)
`define CLP_PV_REG_PCR_ENTRY_14_11                                                                  (32'h1001a8cc)
`define PV_REG_PCR_ENTRY_14_11                                                                      (32'h8cc)
`define CLP_PV_REG_PCR_ENTRY_15_0                                                                   (32'h1001a8d0)
`define PV_REG_PCR_ENTRY_15_0                                                                       (32'h8d0)
`define CLP_PV_REG_PCR_ENTRY_15_1                                                                   (32'h1001a8d4)
`define PV_REG_PCR_ENTRY_15_1                                                                       (32'h8d4)
`define CLP_PV_REG_PCR_ENTRY_15_2                                                                   (32'h1001a8d8)
`define PV_REG_PCR_ENTRY_15_2                                                                       (32'h8d8)
`define CLP_PV_REG_PCR_ENTRY_15_3                                                                   (32'h1001a8dc)
`define PV_REG_PCR_ENTRY_15_3                                                                       (32'h8dc)
`define CLP_PV_REG_PCR_ENTRY_15_4                                                                   (32'h1001a8e0)
`define PV_REG_PCR_ENTRY_15_4                                                                       (32'h8e0)
`define CLP_PV_REG_PCR_ENTRY_15_5                                                                   (32'h1001a8e4)
`define PV_REG_PCR_ENTRY_15_5                                                                       (32'h8e4)
`define CLP_PV_REG_PCR_ENTRY_15_6                                                                   (32'h1001a8e8)
`define PV_REG_PCR_ENTRY_15_6                                                                       (32'h8e8)
`define CLP_PV_REG_PCR_ENTRY_15_7                                                                   (32'h1001a8ec)
`define PV_REG_PCR_ENTRY_15_7                                                                       (32'h8ec)
`define CLP_PV_REG_PCR_ENTRY_15_8                                                                   (32'h1001a8f0)
`define PV_REG_PCR_ENTRY_15_8                                                                       (32'h8f0)
`define CLP_PV_REG_PCR_ENTRY_15_9                                                                   (32'h1001a8f4)
`define PV_REG_PCR_ENTRY_15_9                                                                       (32'h8f4)
`define CLP_PV_REG_PCR_ENTRY_15_10                                                                  (32'h1001a8f8)
`define PV_REG_PCR_ENTRY_15_10                                                                      (32'h8f8)
`define CLP_PV_REG_PCR_ENTRY_15_11                                                                  (32'h1001a8fc)
`define PV_REG_PCR_ENTRY_15_11                                                                      (32'h8fc)
`define CLP_PV_REG_PCR_ENTRY_16_0                                                                   (32'h1001a900)
`define PV_REG_PCR_ENTRY_16_0                                                                       (32'h900)
`define CLP_PV_REG_PCR_ENTRY_16_1                                                                   (32'h1001a904)
`define PV_REG_PCR_ENTRY_16_1                                                                       (32'h904)
`define CLP_PV_REG_PCR_ENTRY_16_2                                                                   (32'h1001a908)
`define PV_REG_PCR_ENTRY_16_2                                                                       (32'h908)
`define CLP_PV_REG_PCR_ENTRY_16_3                                                                   (32'h1001a90c)
`define PV_REG_PCR_ENTRY_16_3                                                                       (32'h90c)
`define CLP_PV_REG_PCR_ENTRY_16_4                                                                   (32'h1001a910)
`define PV_REG_PCR_ENTRY_16_4                                                                       (32'h910)
`define CLP_PV_REG_PCR_ENTRY_16_5                                                                   (32'h1001a914)
`define PV_REG_PCR_ENTRY_16_5                                                                       (32'h914)
`define CLP_PV_REG_PCR_ENTRY_16_6                                                                   (32'h1001a918)
`define PV_REG_PCR_ENTRY_16_6                                                                       (32'h918)
`define CLP_PV_REG_PCR_ENTRY_16_7                                                                   (32'h1001a91c)
`define PV_REG_PCR_ENTRY_16_7                                                                       (32'h91c)
`define CLP_PV_REG_PCR_ENTRY_16_8                                                                   (32'h1001a920)
`define PV_REG_PCR_ENTRY_16_8                                                                       (32'h920)
`define CLP_PV_REG_PCR_ENTRY_16_9                                                                   (32'h1001a924)
`define PV_REG_PCR_ENTRY_16_9                                                                       (32'h924)
`define CLP_PV_REG_PCR_ENTRY_16_10                                                                  (32'h1001a928)
`define PV_REG_PCR_ENTRY_16_10                                                                      (32'h928)
`define CLP_PV_REG_PCR_ENTRY_16_11                                                                  (32'h1001a92c)
`define PV_REG_PCR_ENTRY_16_11                                                                      (32'h92c)
`define CLP_PV_REG_PCR_ENTRY_17_0                                                                   (32'h1001a930)
`define PV_REG_PCR_ENTRY_17_0                                                                       (32'h930)
`define CLP_PV_REG_PCR_ENTRY_17_1                                                                   (32'h1001a934)
`define PV_REG_PCR_ENTRY_17_1                                                                       (32'h934)
`define CLP_PV_REG_PCR_ENTRY_17_2                                                                   (32'h1001a938)
`define PV_REG_PCR_ENTRY_17_2                                                                       (32'h938)
`define CLP_PV_REG_PCR_ENTRY_17_3                                                                   (32'h1001a93c)
`define PV_REG_PCR_ENTRY_17_3                                                                       (32'h93c)
`define CLP_PV_REG_PCR_ENTRY_17_4                                                                   (32'h1001a940)
`define PV_REG_PCR_ENTRY_17_4                                                                       (32'h940)
`define CLP_PV_REG_PCR_ENTRY_17_5                                                                   (32'h1001a944)
`define PV_REG_PCR_ENTRY_17_5                                                                       (32'h944)
`define CLP_PV_REG_PCR_ENTRY_17_6                                                                   (32'h1001a948)
`define PV_REG_PCR_ENTRY_17_6                                                                       (32'h948)
`define CLP_PV_REG_PCR_ENTRY_17_7                                                                   (32'h1001a94c)
`define PV_REG_PCR_ENTRY_17_7                                                                       (32'h94c)
`define CLP_PV_REG_PCR_ENTRY_17_8                                                                   (32'h1001a950)
`define PV_REG_PCR_ENTRY_17_8                                                                       (32'h950)
`define CLP_PV_REG_PCR_ENTRY_17_9                                                                   (32'h1001a954)
`define PV_REG_PCR_ENTRY_17_9                                                                       (32'h954)
`define CLP_PV_REG_PCR_ENTRY_17_10                                                                  (32'h1001a958)
`define PV_REG_PCR_ENTRY_17_10                                                                      (32'h958)
`define CLP_PV_REG_PCR_ENTRY_17_11                                                                  (32'h1001a95c)
`define PV_REG_PCR_ENTRY_17_11                                                                      (32'h95c)
`define CLP_PV_REG_PCR_ENTRY_18_0                                                                   (32'h1001a960)
`define PV_REG_PCR_ENTRY_18_0                                                                       (32'h960)
`define CLP_PV_REG_PCR_ENTRY_18_1                                                                   (32'h1001a964)
`define PV_REG_PCR_ENTRY_18_1                                                                       (32'h964)
`define CLP_PV_REG_PCR_ENTRY_18_2                                                                   (32'h1001a968)
`define PV_REG_PCR_ENTRY_18_2                                                                       (32'h968)
`define CLP_PV_REG_PCR_ENTRY_18_3                                                                   (32'h1001a96c)
`define PV_REG_PCR_ENTRY_18_3                                                                       (32'h96c)
`define CLP_PV_REG_PCR_ENTRY_18_4                                                                   (32'h1001a970)
`define PV_REG_PCR_ENTRY_18_4                                                                       (32'h970)
`define CLP_PV_REG_PCR_ENTRY_18_5                                                                   (32'h1001a974)
`define PV_REG_PCR_ENTRY_18_5                                                                       (32'h974)
`define CLP_PV_REG_PCR_ENTRY_18_6                                                                   (32'h1001a978)
`define PV_REG_PCR_ENTRY_18_6                                                                       (32'h978)
`define CLP_PV_REG_PCR_ENTRY_18_7                                                                   (32'h1001a97c)
`define PV_REG_PCR_ENTRY_18_7                                                                       (32'h97c)
`define CLP_PV_REG_PCR_ENTRY_18_8                                                                   (32'h1001a980)
`define PV_REG_PCR_ENTRY_18_8                                                                       (32'h980)
`define CLP_PV_REG_PCR_ENTRY_18_9                                                                   (32'h1001a984)
`define PV_REG_PCR_ENTRY_18_9                                                                       (32'h984)
`define CLP_PV_REG_PCR_ENTRY_18_10                                                                  (32'h1001a988)
`define PV_REG_PCR_ENTRY_18_10                                                                      (32'h988)
`define CLP_PV_REG_PCR_ENTRY_18_11                                                                  (32'h1001a98c)
`define PV_REG_PCR_ENTRY_18_11                                                                      (32'h98c)
`define CLP_PV_REG_PCR_ENTRY_19_0                                                                   (32'h1001a990)
`define PV_REG_PCR_ENTRY_19_0                                                                       (32'h990)
`define CLP_PV_REG_PCR_ENTRY_19_1                                                                   (32'h1001a994)
`define PV_REG_PCR_ENTRY_19_1                                                                       (32'h994)
`define CLP_PV_REG_PCR_ENTRY_19_2                                                                   (32'h1001a998)
`define PV_REG_PCR_ENTRY_19_2                                                                       (32'h998)
`define CLP_PV_REG_PCR_ENTRY_19_3                                                                   (32'h1001a99c)
`define PV_REG_PCR_ENTRY_19_3                                                                       (32'h99c)
`define CLP_PV_REG_PCR_ENTRY_19_4                                                                   (32'h1001a9a0)
`define PV_REG_PCR_ENTRY_19_4                                                                       (32'h9a0)
`define CLP_PV_REG_PCR_ENTRY_19_5                                                                   (32'h1001a9a4)
`define PV_REG_PCR_ENTRY_19_5                                                                       (32'h9a4)
`define CLP_PV_REG_PCR_ENTRY_19_6                                                                   (32'h1001a9a8)
`define PV_REG_PCR_ENTRY_19_6                                                                       (32'h9a8)
`define CLP_PV_REG_PCR_ENTRY_19_7                                                                   (32'h1001a9ac)
`define PV_REG_PCR_ENTRY_19_7                                                                       (32'h9ac)
`define CLP_PV_REG_PCR_ENTRY_19_8                                                                   (32'h1001a9b0)
`define PV_REG_PCR_ENTRY_19_8                                                                       (32'h9b0)
`define CLP_PV_REG_PCR_ENTRY_19_9                                                                   (32'h1001a9b4)
`define PV_REG_PCR_ENTRY_19_9                                                                       (32'h9b4)
`define CLP_PV_REG_PCR_ENTRY_19_10                                                                  (32'h1001a9b8)
`define PV_REG_PCR_ENTRY_19_10                                                                      (32'h9b8)
`define CLP_PV_REG_PCR_ENTRY_19_11                                                                  (32'h1001a9bc)
`define PV_REG_PCR_ENTRY_19_11                                                                      (32'h9bc)
`define CLP_PV_REG_PCR_ENTRY_20_0                                                                   (32'h1001a9c0)
`define PV_REG_PCR_ENTRY_20_0                                                                       (32'h9c0)
`define CLP_PV_REG_PCR_ENTRY_20_1                                                                   (32'h1001a9c4)
`define PV_REG_PCR_ENTRY_20_1                                                                       (32'h9c4)
`define CLP_PV_REG_PCR_ENTRY_20_2                                                                   (32'h1001a9c8)
`define PV_REG_PCR_ENTRY_20_2                                                                       (32'h9c8)
`define CLP_PV_REG_PCR_ENTRY_20_3                                                                   (32'h1001a9cc)
`define PV_REG_PCR_ENTRY_20_3                                                                       (32'h9cc)
`define CLP_PV_REG_PCR_ENTRY_20_4                                                                   (32'h1001a9d0)
`define PV_REG_PCR_ENTRY_20_4                                                                       (32'h9d0)
`define CLP_PV_REG_PCR_ENTRY_20_5                                                                   (32'h1001a9d4)
`define PV_REG_PCR_ENTRY_20_5                                                                       (32'h9d4)
`define CLP_PV_REG_PCR_ENTRY_20_6                                                                   (32'h1001a9d8)
`define PV_REG_PCR_ENTRY_20_6                                                                       (32'h9d8)
`define CLP_PV_REG_PCR_ENTRY_20_7                                                                   (32'h1001a9dc)
`define PV_REG_PCR_ENTRY_20_7                                                                       (32'h9dc)
`define CLP_PV_REG_PCR_ENTRY_20_8                                                                   (32'h1001a9e0)
`define PV_REG_PCR_ENTRY_20_8                                                                       (32'h9e0)
`define CLP_PV_REG_PCR_ENTRY_20_9                                                                   (32'h1001a9e4)
`define PV_REG_PCR_ENTRY_20_9                                                                       (32'h9e4)
`define CLP_PV_REG_PCR_ENTRY_20_10                                                                  (32'h1001a9e8)
`define PV_REG_PCR_ENTRY_20_10                                                                      (32'h9e8)
`define CLP_PV_REG_PCR_ENTRY_20_11                                                                  (32'h1001a9ec)
`define PV_REG_PCR_ENTRY_20_11                                                                      (32'h9ec)
`define CLP_PV_REG_PCR_ENTRY_21_0                                                                   (32'h1001a9f0)
`define PV_REG_PCR_ENTRY_21_0                                                                       (32'h9f0)
`define CLP_PV_REG_PCR_ENTRY_21_1                                                                   (32'h1001a9f4)
`define PV_REG_PCR_ENTRY_21_1                                                                       (32'h9f4)
`define CLP_PV_REG_PCR_ENTRY_21_2                                                                   (32'h1001a9f8)
`define PV_REG_PCR_ENTRY_21_2                                                                       (32'h9f8)
`define CLP_PV_REG_PCR_ENTRY_21_3                                                                   (32'h1001a9fc)
`define PV_REG_PCR_ENTRY_21_3                                                                       (32'h9fc)
`define CLP_PV_REG_PCR_ENTRY_21_4                                                                   (32'h1001aa00)
`define PV_REG_PCR_ENTRY_21_4                                                                       (32'ha00)
`define CLP_PV_REG_PCR_ENTRY_21_5                                                                   (32'h1001aa04)
`define PV_REG_PCR_ENTRY_21_5                                                                       (32'ha04)
`define CLP_PV_REG_PCR_ENTRY_21_6                                                                   (32'h1001aa08)
`define PV_REG_PCR_ENTRY_21_6                                                                       (32'ha08)
`define CLP_PV_REG_PCR_ENTRY_21_7                                                                   (32'h1001aa0c)
`define PV_REG_PCR_ENTRY_21_7                                                                       (32'ha0c)
`define CLP_PV_REG_PCR_ENTRY_21_8                                                                   (32'h1001aa10)
`define PV_REG_PCR_ENTRY_21_8                                                                       (32'ha10)
`define CLP_PV_REG_PCR_ENTRY_21_9                                                                   (32'h1001aa14)
`define PV_REG_PCR_ENTRY_21_9                                                                       (32'ha14)
`define CLP_PV_REG_PCR_ENTRY_21_10                                                                  (32'h1001aa18)
`define PV_REG_PCR_ENTRY_21_10                                                                      (32'ha18)
`define CLP_PV_REG_PCR_ENTRY_21_11                                                                  (32'h1001aa1c)
`define PV_REG_PCR_ENTRY_21_11                                                                      (32'ha1c)
`define CLP_PV_REG_PCR_ENTRY_22_0                                                                   (32'h1001aa20)
`define PV_REG_PCR_ENTRY_22_0                                                                       (32'ha20)
`define CLP_PV_REG_PCR_ENTRY_22_1                                                                   (32'h1001aa24)
`define PV_REG_PCR_ENTRY_22_1                                                                       (32'ha24)
`define CLP_PV_REG_PCR_ENTRY_22_2                                                                   (32'h1001aa28)
`define PV_REG_PCR_ENTRY_22_2                                                                       (32'ha28)
`define CLP_PV_REG_PCR_ENTRY_22_3                                                                   (32'h1001aa2c)
`define PV_REG_PCR_ENTRY_22_3                                                                       (32'ha2c)
`define CLP_PV_REG_PCR_ENTRY_22_4                                                                   (32'h1001aa30)
`define PV_REG_PCR_ENTRY_22_4                                                                       (32'ha30)
`define CLP_PV_REG_PCR_ENTRY_22_5                                                                   (32'h1001aa34)
`define PV_REG_PCR_ENTRY_22_5                                                                       (32'ha34)
`define CLP_PV_REG_PCR_ENTRY_22_6                                                                   (32'h1001aa38)
`define PV_REG_PCR_ENTRY_22_6                                                                       (32'ha38)
`define CLP_PV_REG_PCR_ENTRY_22_7                                                                   (32'h1001aa3c)
`define PV_REG_PCR_ENTRY_22_7                                                                       (32'ha3c)
`define CLP_PV_REG_PCR_ENTRY_22_8                                                                   (32'h1001aa40)
`define PV_REG_PCR_ENTRY_22_8                                                                       (32'ha40)
`define CLP_PV_REG_PCR_ENTRY_22_9                                                                   (32'h1001aa44)
`define PV_REG_PCR_ENTRY_22_9                                                                       (32'ha44)
`define CLP_PV_REG_PCR_ENTRY_22_10                                                                  (32'h1001aa48)
`define PV_REG_PCR_ENTRY_22_10                                                                      (32'ha48)
`define CLP_PV_REG_PCR_ENTRY_22_11                                                                  (32'h1001aa4c)
`define PV_REG_PCR_ENTRY_22_11                                                                      (32'ha4c)
`define CLP_PV_REG_PCR_ENTRY_23_0                                                                   (32'h1001aa50)
`define PV_REG_PCR_ENTRY_23_0                                                                       (32'ha50)
`define CLP_PV_REG_PCR_ENTRY_23_1                                                                   (32'h1001aa54)
`define PV_REG_PCR_ENTRY_23_1                                                                       (32'ha54)
`define CLP_PV_REG_PCR_ENTRY_23_2                                                                   (32'h1001aa58)
`define PV_REG_PCR_ENTRY_23_2                                                                       (32'ha58)
`define CLP_PV_REG_PCR_ENTRY_23_3                                                                   (32'h1001aa5c)
`define PV_REG_PCR_ENTRY_23_3                                                                       (32'ha5c)
`define CLP_PV_REG_PCR_ENTRY_23_4                                                                   (32'h1001aa60)
`define PV_REG_PCR_ENTRY_23_4                                                                       (32'ha60)
`define CLP_PV_REG_PCR_ENTRY_23_5                                                                   (32'h1001aa64)
`define PV_REG_PCR_ENTRY_23_5                                                                       (32'ha64)
`define CLP_PV_REG_PCR_ENTRY_23_6                                                                   (32'h1001aa68)
`define PV_REG_PCR_ENTRY_23_6                                                                       (32'ha68)
`define CLP_PV_REG_PCR_ENTRY_23_7                                                                   (32'h1001aa6c)
`define PV_REG_PCR_ENTRY_23_7                                                                       (32'ha6c)
`define CLP_PV_REG_PCR_ENTRY_23_8                                                                   (32'h1001aa70)
`define PV_REG_PCR_ENTRY_23_8                                                                       (32'ha70)
`define CLP_PV_REG_PCR_ENTRY_23_9                                                                   (32'h1001aa74)
`define PV_REG_PCR_ENTRY_23_9                                                                       (32'ha74)
`define CLP_PV_REG_PCR_ENTRY_23_10                                                                  (32'h1001aa78)
`define PV_REG_PCR_ENTRY_23_10                                                                      (32'ha78)
`define CLP_PV_REG_PCR_ENTRY_23_11                                                                  (32'h1001aa7c)
`define PV_REG_PCR_ENTRY_23_11                                                                      (32'ha7c)
`define CLP_PV_REG_PCR_ENTRY_24_0                                                                   (32'h1001aa80)
`define PV_REG_PCR_ENTRY_24_0                                                                       (32'ha80)
`define CLP_PV_REG_PCR_ENTRY_24_1                                                                   (32'h1001aa84)
`define PV_REG_PCR_ENTRY_24_1                                                                       (32'ha84)
`define CLP_PV_REG_PCR_ENTRY_24_2                                                                   (32'h1001aa88)
`define PV_REG_PCR_ENTRY_24_2                                                                       (32'ha88)
`define CLP_PV_REG_PCR_ENTRY_24_3                                                                   (32'h1001aa8c)
`define PV_REG_PCR_ENTRY_24_3                                                                       (32'ha8c)
`define CLP_PV_REG_PCR_ENTRY_24_4                                                                   (32'h1001aa90)
`define PV_REG_PCR_ENTRY_24_4                                                                       (32'ha90)
`define CLP_PV_REG_PCR_ENTRY_24_5                                                                   (32'h1001aa94)
`define PV_REG_PCR_ENTRY_24_5                                                                       (32'ha94)
`define CLP_PV_REG_PCR_ENTRY_24_6                                                                   (32'h1001aa98)
`define PV_REG_PCR_ENTRY_24_6                                                                       (32'ha98)
`define CLP_PV_REG_PCR_ENTRY_24_7                                                                   (32'h1001aa9c)
`define PV_REG_PCR_ENTRY_24_7                                                                       (32'ha9c)
`define CLP_PV_REG_PCR_ENTRY_24_8                                                                   (32'h1001aaa0)
`define PV_REG_PCR_ENTRY_24_8                                                                       (32'haa0)
`define CLP_PV_REG_PCR_ENTRY_24_9                                                                   (32'h1001aaa4)
`define PV_REG_PCR_ENTRY_24_9                                                                       (32'haa4)
`define CLP_PV_REG_PCR_ENTRY_24_10                                                                  (32'h1001aaa8)
`define PV_REG_PCR_ENTRY_24_10                                                                      (32'haa8)
`define CLP_PV_REG_PCR_ENTRY_24_11                                                                  (32'h1001aaac)
`define PV_REG_PCR_ENTRY_24_11                                                                      (32'haac)
`define CLP_PV_REG_PCR_ENTRY_25_0                                                                   (32'h1001aab0)
`define PV_REG_PCR_ENTRY_25_0                                                                       (32'hab0)
`define CLP_PV_REG_PCR_ENTRY_25_1                                                                   (32'h1001aab4)
`define PV_REG_PCR_ENTRY_25_1                                                                       (32'hab4)
`define CLP_PV_REG_PCR_ENTRY_25_2                                                                   (32'h1001aab8)
`define PV_REG_PCR_ENTRY_25_2                                                                       (32'hab8)
`define CLP_PV_REG_PCR_ENTRY_25_3                                                                   (32'h1001aabc)
`define PV_REG_PCR_ENTRY_25_3                                                                       (32'habc)
`define CLP_PV_REG_PCR_ENTRY_25_4                                                                   (32'h1001aac0)
`define PV_REG_PCR_ENTRY_25_4                                                                       (32'hac0)
`define CLP_PV_REG_PCR_ENTRY_25_5                                                                   (32'h1001aac4)
`define PV_REG_PCR_ENTRY_25_5                                                                       (32'hac4)
`define CLP_PV_REG_PCR_ENTRY_25_6                                                                   (32'h1001aac8)
`define PV_REG_PCR_ENTRY_25_6                                                                       (32'hac8)
`define CLP_PV_REG_PCR_ENTRY_25_7                                                                   (32'h1001aacc)
`define PV_REG_PCR_ENTRY_25_7                                                                       (32'hacc)
`define CLP_PV_REG_PCR_ENTRY_25_8                                                                   (32'h1001aad0)
`define PV_REG_PCR_ENTRY_25_8                                                                       (32'had0)
`define CLP_PV_REG_PCR_ENTRY_25_9                                                                   (32'h1001aad4)
`define PV_REG_PCR_ENTRY_25_9                                                                       (32'had4)
`define CLP_PV_REG_PCR_ENTRY_25_10                                                                  (32'h1001aad8)
`define PV_REG_PCR_ENTRY_25_10                                                                      (32'had8)
`define CLP_PV_REG_PCR_ENTRY_25_11                                                                  (32'h1001aadc)
`define PV_REG_PCR_ENTRY_25_11                                                                      (32'hadc)
`define CLP_PV_REG_PCR_ENTRY_26_0                                                                   (32'h1001aae0)
`define PV_REG_PCR_ENTRY_26_0                                                                       (32'hae0)
`define CLP_PV_REG_PCR_ENTRY_26_1                                                                   (32'h1001aae4)
`define PV_REG_PCR_ENTRY_26_1                                                                       (32'hae4)
`define CLP_PV_REG_PCR_ENTRY_26_2                                                                   (32'h1001aae8)
`define PV_REG_PCR_ENTRY_26_2                                                                       (32'hae8)
`define CLP_PV_REG_PCR_ENTRY_26_3                                                                   (32'h1001aaec)
`define PV_REG_PCR_ENTRY_26_3                                                                       (32'haec)
`define CLP_PV_REG_PCR_ENTRY_26_4                                                                   (32'h1001aaf0)
`define PV_REG_PCR_ENTRY_26_4                                                                       (32'haf0)
`define CLP_PV_REG_PCR_ENTRY_26_5                                                                   (32'h1001aaf4)
`define PV_REG_PCR_ENTRY_26_5                                                                       (32'haf4)
`define CLP_PV_REG_PCR_ENTRY_26_6                                                                   (32'h1001aaf8)
`define PV_REG_PCR_ENTRY_26_6                                                                       (32'haf8)
`define CLP_PV_REG_PCR_ENTRY_26_7                                                                   (32'h1001aafc)
`define PV_REG_PCR_ENTRY_26_7                                                                       (32'hafc)
`define CLP_PV_REG_PCR_ENTRY_26_8                                                                   (32'h1001ab00)
`define PV_REG_PCR_ENTRY_26_8                                                                       (32'hb00)
`define CLP_PV_REG_PCR_ENTRY_26_9                                                                   (32'h1001ab04)
`define PV_REG_PCR_ENTRY_26_9                                                                       (32'hb04)
`define CLP_PV_REG_PCR_ENTRY_26_10                                                                  (32'h1001ab08)
`define PV_REG_PCR_ENTRY_26_10                                                                      (32'hb08)
`define CLP_PV_REG_PCR_ENTRY_26_11                                                                  (32'h1001ab0c)
`define PV_REG_PCR_ENTRY_26_11                                                                      (32'hb0c)
`define CLP_PV_REG_PCR_ENTRY_27_0                                                                   (32'h1001ab10)
`define PV_REG_PCR_ENTRY_27_0                                                                       (32'hb10)
`define CLP_PV_REG_PCR_ENTRY_27_1                                                                   (32'h1001ab14)
`define PV_REG_PCR_ENTRY_27_1                                                                       (32'hb14)
`define CLP_PV_REG_PCR_ENTRY_27_2                                                                   (32'h1001ab18)
`define PV_REG_PCR_ENTRY_27_2                                                                       (32'hb18)
`define CLP_PV_REG_PCR_ENTRY_27_3                                                                   (32'h1001ab1c)
`define PV_REG_PCR_ENTRY_27_3                                                                       (32'hb1c)
`define CLP_PV_REG_PCR_ENTRY_27_4                                                                   (32'h1001ab20)
`define PV_REG_PCR_ENTRY_27_4                                                                       (32'hb20)
`define CLP_PV_REG_PCR_ENTRY_27_5                                                                   (32'h1001ab24)
`define PV_REG_PCR_ENTRY_27_5                                                                       (32'hb24)
`define CLP_PV_REG_PCR_ENTRY_27_6                                                                   (32'h1001ab28)
`define PV_REG_PCR_ENTRY_27_6                                                                       (32'hb28)
`define CLP_PV_REG_PCR_ENTRY_27_7                                                                   (32'h1001ab2c)
`define PV_REG_PCR_ENTRY_27_7                                                                       (32'hb2c)
`define CLP_PV_REG_PCR_ENTRY_27_8                                                                   (32'h1001ab30)
`define PV_REG_PCR_ENTRY_27_8                                                                       (32'hb30)
`define CLP_PV_REG_PCR_ENTRY_27_9                                                                   (32'h1001ab34)
`define PV_REG_PCR_ENTRY_27_9                                                                       (32'hb34)
`define CLP_PV_REG_PCR_ENTRY_27_10                                                                  (32'h1001ab38)
`define PV_REG_PCR_ENTRY_27_10                                                                      (32'hb38)
`define CLP_PV_REG_PCR_ENTRY_27_11                                                                  (32'h1001ab3c)
`define PV_REG_PCR_ENTRY_27_11                                                                      (32'hb3c)
`define CLP_PV_REG_PCR_ENTRY_28_0                                                                   (32'h1001ab40)
`define PV_REG_PCR_ENTRY_28_0                                                                       (32'hb40)
`define CLP_PV_REG_PCR_ENTRY_28_1                                                                   (32'h1001ab44)
`define PV_REG_PCR_ENTRY_28_1                                                                       (32'hb44)
`define CLP_PV_REG_PCR_ENTRY_28_2                                                                   (32'h1001ab48)
`define PV_REG_PCR_ENTRY_28_2                                                                       (32'hb48)
`define CLP_PV_REG_PCR_ENTRY_28_3                                                                   (32'h1001ab4c)
`define PV_REG_PCR_ENTRY_28_3                                                                       (32'hb4c)
`define CLP_PV_REG_PCR_ENTRY_28_4                                                                   (32'h1001ab50)
`define PV_REG_PCR_ENTRY_28_4                                                                       (32'hb50)
`define CLP_PV_REG_PCR_ENTRY_28_5                                                                   (32'h1001ab54)
`define PV_REG_PCR_ENTRY_28_5                                                                       (32'hb54)
`define CLP_PV_REG_PCR_ENTRY_28_6                                                                   (32'h1001ab58)
`define PV_REG_PCR_ENTRY_28_6                                                                       (32'hb58)
`define CLP_PV_REG_PCR_ENTRY_28_7                                                                   (32'h1001ab5c)
`define PV_REG_PCR_ENTRY_28_7                                                                       (32'hb5c)
`define CLP_PV_REG_PCR_ENTRY_28_8                                                                   (32'h1001ab60)
`define PV_REG_PCR_ENTRY_28_8                                                                       (32'hb60)
`define CLP_PV_REG_PCR_ENTRY_28_9                                                                   (32'h1001ab64)
`define PV_REG_PCR_ENTRY_28_9                                                                       (32'hb64)
`define CLP_PV_REG_PCR_ENTRY_28_10                                                                  (32'h1001ab68)
`define PV_REG_PCR_ENTRY_28_10                                                                      (32'hb68)
`define CLP_PV_REG_PCR_ENTRY_28_11                                                                  (32'h1001ab6c)
`define PV_REG_PCR_ENTRY_28_11                                                                      (32'hb6c)
`define CLP_PV_REG_PCR_ENTRY_29_0                                                                   (32'h1001ab70)
`define PV_REG_PCR_ENTRY_29_0                                                                       (32'hb70)
`define CLP_PV_REG_PCR_ENTRY_29_1                                                                   (32'h1001ab74)
`define PV_REG_PCR_ENTRY_29_1                                                                       (32'hb74)
`define CLP_PV_REG_PCR_ENTRY_29_2                                                                   (32'h1001ab78)
`define PV_REG_PCR_ENTRY_29_2                                                                       (32'hb78)
`define CLP_PV_REG_PCR_ENTRY_29_3                                                                   (32'h1001ab7c)
`define PV_REG_PCR_ENTRY_29_3                                                                       (32'hb7c)
`define CLP_PV_REG_PCR_ENTRY_29_4                                                                   (32'h1001ab80)
`define PV_REG_PCR_ENTRY_29_4                                                                       (32'hb80)
`define CLP_PV_REG_PCR_ENTRY_29_5                                                                   (32'h1001ab84)
`define PV_REG_PCR_ENTRY_29_5                                                                       (32'hb84)
`define CLP_PV_REG_PCR_ENTRY_29_6                                                                   (32'h1001ab88)
`define PV_REG_PCR_ENTRY_29_6                                                                       (32'hb88)
`define CLP_PV_REG_PCR_ENTRY_29_7                                                                   (32'h1001ab8c)
`define PV_REG_PCR_ENTRY_29_7                                                                       (32'hb8c)
`define CLP_PV_REG_PCR_ENTRY_29_8                                                                   (32'h1001ab90)
`define PV_REG_PCR_ENTRY_29_8                                                                       (32'hb90)
`define CLP_PV_REG_PCR_ENTRY_29_9                                                                   (32'h1001ab94)
`define PV_REG_PCR_ENTRY_29_9                                                                       (32'hb94)
`define CLP_PV_REG_PCR_ENTRY_29_10                                                                  (32'h1001ab98)
`define PV_REG_PCR_ENTRY_29_10                                                                      (32'hb98)
`define CLP_PV_REG_PCR_ENTRY_29_11                                                                  (32'h1001ab9c)
`define PV_REG_PCR_ENTRY_29_11                                                                      (32'hb9c)
`define CLP_PV_REG_PCR_ENTRY_30_0                                                                   (32'h1001aba0)
`define PV_REG_PCR_ENTRY_30_0                                                                       (32'hba0)
`define CLP_PV_REG_PCR_ENTRY_30_1                                                                   (32'h1001aba4)
`define PV_REG_PCR_ENTRY_30_1                                                                       (32'hba4)
`define CLP_PV_REG_PCR_ENTRY_30_2                                                                   (32'h1001aba8)
`define PV_REG_PCR_ENTRY_30_2                                                                       (32'hba8)
`define CLP_PV_REG_PCR_ENTRY_30_3                                                                   (32'h1001abac)
`define PV_REG_PCR_ENTRY_30_3                                                                       (32'hbac)
`define CLP_PV_REG_PCR_ENTRY_30_4                                                                   (32'h1001abb0)
`define PV_REG_PCR_ENTRY_30_4                                                                       (32'hbb0)
`define CLP_PV_REG_PCR_ENTRY_30_5                                                                   (32'h1001abb4)
`define PV_REG_PCR_ENTRY_30_5                                                                       (32'hbb4)
`define CLP_PV_REG_PCR_ENTRY_30_6                                                                   (32'h1001abb8)
`define PV_REG_PCR_ENTRY_30_6                                                                       (32'hbb8)
`define CLP_PV_REG_PCR_ENTRY_30_7                                                                   (32'h1001abbc)
`define PV_REG_PCR_ENTRY_30_7                                                                       (32'hbbc)
`define CLP_PV_REG_PCR_ENTRY_30_8                                                                   (32'h1001abc0)
`define PV_REG_PCR_ENTRY_30_8                                                                       (32'hbc0)
`define CLP_PV_REG_PCR_ENTRY_30_9                                                                   (32'h1001abc4)
`define PV_REG_PCR_ENTRY_30_9                                                                       (32'hbc4)
`define CLP_PV_REG_PCR_ENTRY_30_10                                                                  (32'h1001abc8)
`define PV_REG_PCR_ENTRY_30_10                                                                      (32'hbc8)
`define CLP_PV_REG_PCR_ENTRY_30_11                                                                  (32'h1001abcc)
`define PV_REG_PCR_ENTRY_30_11                                                                      (32'hbcc)
`define CLP_PV_REG_PCR_ENTRY_31_0                                                                   (32'h1001abd0)
`define PV_REG_PCR_ENTRY_31_0                                                                       (32'hbd0)
`define CLP_PV_REG_PCR_ENTRY_31_1                                                                   (32'h1001abd4)
`define PV_REG_PCR_ENTRY_31_1                                                                       (32'hbd4)
`define CLP_PV_REG_PCR_ENTRY_31_2                                                                   (32'h1001abd8)
`define PV_REG_PCR_ENTRY_31_2                                                                       (32'hbd8)
`define CLP_PV_REG_PCR_ENTRY_31_3                                                                   (32'h1001abdc)
`define PV_REG_PCR_ENTRY_31_3                                                                       (32'hbdc)
`define CLP_PV_REG_PCR_ENTRY_31_4                                                                   (32'h1001abe0)
`define PV_REG_PCR_ENTRY_31_4                                                                       (32'hbe0)
`define CLP_PV_REG_PCR_ENTRY_31_5                                                                   (32'h1001abe4)
`define PV_REG_PCR_ENTRY_31_5                                                                       (32'hbe4)
`define CLP_PV_REG_PCR_ENTRY_31_6                                                                   (32'h1001abe8)
`define PV_REG_PCR_ENTRY_31_6                                                                       (32'hbe8)
`define CLP_PV_REG_PCR_ENTRY_31_7                                                                   (32'h1001abec)
`define PV_REG_PCR_ENTRY_31_7                                                                       (32'hbec)
`define CLP_PV_REG_PCR_ENTRY_31_8                                                                   (32'h1001abf0)
`define PV_REG_PCR_ENTRY_31_8                                                                       (32'hbf0)
`define CLP_PV_REG_PCR_ENTRY_31_9                                                                   (32'h1001abf4)
`define PV_REG_PCR_ENTRY_31_9                                                                       (32'hbf4)
`define CLP_PV_REG_PCR_ENTRY_31_10                                                                  (32'h1001abf8)
`define PV_REG_PCR_ENTRY_31_10                                                                      (32'hbf8)
`define CLP_PV_REG_PCR_ENTRY_31_11                                                                  (32'h1001abfc)
`define PV_REG_PCR_ENTRY_31_11                                                                      (32'hbfc)
`define CLP_DV_REG_BASE_ADDR                                                                        (32'h1001c000)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_0                                                            (32'h1001c000)
`define DV_REG_STICKYDATAVAULTCTRL_0                                                                (32'h0)
`define DV_REG_STICKYDATAVAULTCTRL_0_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_0_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_1                                                            (32'h1001c004)
`define DV_REG_STICKYDATAVAULTCTRL_1                                                                (32'h4)
`define DV_REG_STICKYDATAVAULTCTRL_1_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_1_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_2                                                            (32'h1001c008)
`define DV_REG_STICKYDATAVAULTCTRL_2                                                                (32'h8)
`define DV_REG_STICKYDATAVAULTCTRL_2_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_2_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_3                                                            (32'h1001c00c)
`define DV_REG_STICKYDATAVAULTCTRL_3                                                                (32'hc)
`define DV_REG_STICKYDATAVAULTCTRL_3_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_3_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_4                                                            (32'h1001c010)
`define DV_REG_STICKYDATAVAULTCTRL_4                                                                (32'h10)
`define DV_REG_STICKYDATAVAULTCTRL_4_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_4_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_5                                                            (32'h1001c014)
`define DV_REG_STICKYDATAVAULTCTRL_5                                                                (32'h14)
`define DV_REG_STICKYDATAVAULTCTRL_5_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_5_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_6                                                            (32'h1001c018)
`define DV_REG_STICKYDATAVAULTCTRL_6                                                                (32'h18)
`define DV_REG_STICKYDATAVAULTCTRL_6_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_6_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_7                                                            (32'h1001c01c)
`define DV_REG_STICKYDATAVAULTCTRL_7                                                                (32'h1c)
`define DV_REG_STICKYDATAVAULTCTRL_7_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_7_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_8                                                            (32'h1001c020)
`define DV_REG_STICKYDATAVAULTCTRL_8                                                                (32'h20)
`define DV_REG_STICKYDATAVAULTCTRL_8_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_8_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKYDATAVAULTCTRL_9                                                            (32'h1001c024)
`define DV_REG_STICKYDATAVAULTCTRL_9                                                                (32'h24)
`define DV_REG_STICKYDATAVAULTCTRL_9_LOCK_ENTRY_LOW                                                 (0)
`define DV_REG_STICKYDATAVAULTCTRL_9_LOCK_ENTRY_MASK                                                (32'h1)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_0                                                      (32'h1001c028)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_0                                                          (32'h28)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_1                                                      (32'h1001c02c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_1                                                          (32'h2c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_2                                                      (32'h1001c030)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_2                                                          (32'h30)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_3                                                      (32'h1001c034)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_3                                                          (32'h34)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_4                                                      (32'h1001c038)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_4                                                          (32'h38)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_5                                                      (32'h1001c03c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_5                                                          (32'h3c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_6                                                      (32'h1001c040)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_6                                                          (32'h40)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_7                                                      (32'h1001c044)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_7                                                          (32'h44)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_8                                                      (32'h1001c048)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_8                                                          (32'h48)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_9                                                      (32'h1001c04c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_9                                                          (32'h4c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_10                                                     (32'h1001c050)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_10                                                         (32'h50)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_0_11                                                     (32'h1001c054)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_0_11                                                         (32'h54)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_0                                                      (32'h1001c058)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_0                                                          (32'h58)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_1                                                      (32'h1001c05c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_1                                                          (32'h5c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_2                                                      (32'h1001c060)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_2                                                          (32'h60)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_3                                                      (32'h1001c064)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_3                                                          (32'h64)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_4                                                      (32'h1001c068)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_4                                                          (32'h68)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_5                                                      (32'h1001c06c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_5                                                          (32'h6c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_6                                                      (32'h1001c070)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_6                                                          (32'h70)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_7                                                      (32'h1001c074)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_7                                                          (32'h74)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_8                                                      (32'h1001c078)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_8                                                          (32'h78)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_9                                                      (32'h1001c07c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_9                                                          (32'h7c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_10                                                     (32'h1001c080)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_10                                                         (32'h80)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_1_11                                                     (32'h1001c084)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_1_11                                                         (32'h84)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_0                                                      (32'h1001c088)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_0                                                          (32'h88)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_1                                                      (32'h1001c08c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_1                                                          (32'h8c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_2                                                      (32'h1001c090)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_2                                                          (32'h90)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_3                                                      (32'h1001c094)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_3                                                          (32'h94)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_4                                                      (32'h1001c098)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_4                                                          (32'h98)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_5                                                      (32'h1001c09c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_5                                                          (32'h9c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_6                                                      (32'h1001c0a0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_6                                                          (32'ha0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_7                                                      (32'h1001c0a4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_7                                                          (32'ha4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_8                                                      (32'h1001c0a8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_8                                                          (32'ha8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_9                                                      (32'h1001c0ac)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_9                                                          (32'hac)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_10                                                     (32'h1001c0b0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_10                                                         (32'hb0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_2_11                                                     (32'h1001c0b4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_2_11                                                         (32'hb4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_0                                                      (32'h1001c0b8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_0                                                          (32'hb8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_1                                                      (32'h1001c0bc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_1                                                          (32'hbc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_2                                                      (32'h1001c0c0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_2                                                          (32'hc0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_3                                                      (32'h1001c0c4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_3                                                          (32'hc4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_4                                                      (32'h1001c0c8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_4                                                          (32'hc8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_5                                                      (32'h1001c0cc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_5                                                          (32'hcc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_6                                                      (32'h1001c0d0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_6                                                          (32'hd0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_7                                                      (32'h1001c0d4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_7                                                          (32'hd4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_8                                                      (32'h1001c0d8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_8                                                          (32'hd8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_9                                                      (32'h1001c0dc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_9                                                          (32'hdc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_10                                                     (32'h1001c0e0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_10                                                         (32'he0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_3_11                                                     (32'h1001c0e4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_3_11                                                         (32'he4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_0                                                      (32'h1001c0e8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_0                                                          (32'he8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_1                                                      (32'h1001c0ec)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_1                                                          (32'hec)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_2                                                      (32'h1001c0f0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_2                                                          (32'hf0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_3                                                      (32'h1001c0f4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_3                                                          (32'hf4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_4                                                      (32'h1001c0f8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_4                                                          (32'hf8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_5                                                      (32'h1001c0fc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_5                                                          (32'hfc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_6                                                      (32'h1001c100)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_6                                                          (32'h100)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_7                                                      (32'h1001c104)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_7                                                          (32'h104)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_8                                                      (32'h1001c108)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_8                                                          (32'h108)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_9                                                      (32'h1001c10c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_9                                                          (32'h10c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_10                                                     (32'h1001c110)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_10                                                         (32'h110)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_4_11                                                     (32'h1001c114)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_4_11                                                         (32'h114)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_0                                                      (32'h1001c118)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_0                                                          (32'h118)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_1                                                      (32'h1001c11c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_1                                                          (32'h11c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_2                                                      (32'h1001c120)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_2                                                          (32'h120)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_3                                                      (32'h1001c124)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_3                                                          (32'h124)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_4                                                      (32'h1001c128)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_4                                                          (32'h128)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_5                                                      (32'h1001c12c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_5                                                          (32'h12c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_6                                                      (32'h1001c130)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_6                                                          (32'h130)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_7                                                      (32'h1001c134)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_7                                                          (32'h134)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_8                                                      (32'h1001c138)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_8                                                          (32'h138)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_9                                                      (32'h1001c13c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_9                                                          (32'h13c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_10                                                     (32'h1001c140)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_10                                                         (32'h140)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_5_11                                                     (32'h1001c144)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_5_11                                                         (32'h144)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_0                                                      (32'h1001c148)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_0                                                          (32'h148)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_1                                                      (32'h1001c14c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_1                                                          (32'h14c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_2                                                      (32'h1001c150)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_2                                                          (32'h150)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_3                                                      (32'h1001c154)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_3                                                          (32'h154)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_4                                                      (32'h1001c158)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_4                                                          (32'h158)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_5                                                      (32'h1001c15c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_5                                                          (32'h15c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_6                                                      (32'h1001c160)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_6                                                          (32'h160)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_7                                                      (32'h1001c164)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_7                                                          (32'h164)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_8                                                      (32'h1001c168)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_8                                                          (32'h168)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_9                                                      (32'h1001c16c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_9                                                          (32'h16c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_10                                                     (32'h1001c170)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_10                                                         (32'h170)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_6_11                                                     (32'h1001c174)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_6_11                                                         (32'h174)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_0                                                      (32'h1001c178)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_0                                                          (32'h178)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_1                                                      (32'h1001c17c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_1                                                          (32'h17c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_2                                                      (32'h1001c180)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_2                                                          (32'h180)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_3                                                      (32'h1001c184)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_3                                                          (32'h184)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_4                                                      (32'h1001c188)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_4                                                          (32'h188)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_5                                                      (32'h1001c18c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_5                                                          (32'h18c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_6                                                      (32'h1001c190)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_6                                                          (32'h190)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_7                                                      (32'h1001c194)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_7                                                          (32'h194)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_8                                                      (32'h1001c198)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_8                                                          (32'h198)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_9                                                      (32'h1001c19c)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_9                                                          (32'h19c)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_10                                                     (32'h1001c1a0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_10                                                         (32'h1a0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_7_11                                                     (32'h1001c1a4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_7_11                                                         (32'h1a4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_0                                                      (32'h1001c1a8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_0                                                          (32'h1a8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_1                                                      (32'h1001c1ac)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_1                                                          (32'h1ac)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_2                                                      (32'h1001c1b0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_2                                                          (32'h1b0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_3                                                      (32'h1001c1b4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_3                                                          (32'h1b4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_4                                                      (32'h1001c1b8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_4                                                          (32'h1b8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_5                                                      (32'h1001c1bc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_5                                                          (32'h1bc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_6                                                      (32'h1001c1c0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_6                                                          (32'h1c0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_7                                                      (32'h1001c1c4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_7                                                          (32'h1c4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_8                                                      (32'h1001c1c8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_8                                                          (32'h1c8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_9                                                      (32'h1001c1cc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_9                                                          (32'h1cc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_10                                                     (32'h1001c1d0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_10                                                         (32'h1d0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_8_11                                                     (32'h1001c1d4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_8_11                                                         (32'h1d4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_0                                                      (32'h1001c1d8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_0                                                          (32'h1d8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_1                                                      (32'h1001c1dc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_1                                                          (32'h1dc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_2                                                      (32'h1001c1e0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_2                                                          (32'h1e0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_3                                                      (32'h1001c1e4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_3                                                          (32'h1e4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_4                                                      (32'h1001c1e8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_4                                                          (32'h1e8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_5                                                      (32'h1001c1ec)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_5                                                          (32'h1ec)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_6                                                      (32'h1001c1f0)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_6                                                          (32'h1f0)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_7                                                      (32'h1001c1f4)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_7                                                          (32'h1f4)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_8                                                      (32'h1001c1f8)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_8                                                          (32'h1f8)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_9                                                      (32'h1001c1fc)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_9                                                          (32'h1fc)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_10                                                     (32'h1001c200)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_10                                                         (32'h200)
`define CLP_DV_REG_STICKY_DATA_VAULT_ENTRY_9_11                                                     (32'h1001c204)
`define DV_REG_STICKY_DATA_VAULT_ENTRY_9_11                                                         (32'h204)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_0                                                         (32'h1001c208)
`define DV_REG_NONSTICKYDATAVAULTCTRL_0                                                             (32'h208)
`define DV_REG_NONSTICKYDATAVAULTCTRL_0_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_0_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_1                                                         (32'h1001c20c)
`define DV_REG_NONSTICKYDATAVAULTCTRL_1                                                             (32'h20c)
`define DV_REG_NONSTICKYDATAVAULTCTRL_1_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_1_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_2                                                         (32'h1001c210)
`define DV_REG_NONSTICKYDATAVAULTCTRL_2                                                             (32'h210)
`define DV_REG_NONSTICKYDATAVAULTCTRL_2_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_2_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_3                                                         (32'h1001c214)
`define DV_REG_NONSTICKYDATAVAULTCTRL_3                                                             (32'h214)
`define DV_REG_NONSTICKYDATAVAULTCTRL_3_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_3_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_4                                                         (32'h1001c218)
`define DV_REG_NONSTICKYDATAVAULTCTRL_4                                                             (32'h218)
`define DV_REG_NONSTICKYDATAVAULTCTRL_4_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_4_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_5                                                         (32'h1001c21c)
`define DV_REG_NONSTICKYDATAVAULTCTRL_5                                                             (32'h21c)
`define DV_REG_NONSTICKYDATAVAULTCTRL_5_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_5_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_6                                                         (32'h1001c220)
`define DV_REG_NONSTICKYDATAVAULTCTRL_6                                                             (32'h220)
`define DV_REG_NONSTICKYDATAVAULTCTRL_6_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_6_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_7                                                         (32'h1001c224)
`define DV_REG_NONSTICKYDATAVAULTCTRL_7                                                             (32'h224)
`define DV_REG_NONSTICKYDATAVAULTCTRL_7_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_7_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_8                                                         (32'h1001c228)
`define DV_REG_NONSTICKYDATAVAULTCTRL_8                                                             (32'h228)
`define DV_REG_NONSTICKYDATAVAULTCTRL_8_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_8_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKYDATAVAULTCTRL_9                                                         (32'h1001c22c)
`define DV_REG_NONSTICKYDATAVAULTCTRL_9                                                             (32'h22c)
`define DV_REG_NONSTICKYDATAVAULTCTRL_9_LOCK_ENTRY_LOW                                              (0)
`define DV_REG_NONSTICKYDATAVAULTCTRL_9_LOCK_ENTRY_MASK                                             (32'h1)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_0                                                   (32'h1001c230)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_0                                                       (32'h230)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_1                                                   (32'h1001c234)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_1                                                       (32'h234)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_2                                                   (32'h1001c238)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_2                                                       (32'h238)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_3                                                   (32'h1001c23c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_3                                                       (32'h23c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_4                                                   (32'h1001c240)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_4                                                       (32'h240)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_5                                                   (32'h1001c244)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_5                                                       (32'h244)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_6                                                   (32'h1001c248)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_6                                                       (32'h248)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_7                                                   (32'h1001c24c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_7                                                       (32'h24c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_8                                                   (32'h1001c250)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_8                                                       (32'h250)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_9                                                   (32'h1001c254)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_9                                                       (32'h254)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_10                                                  (32'h1001c258)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_10                                                      (32'h258)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_11                                                  (32'h1001c25c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_0_11                                                      (32'h25c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_0                                                   (32'h1001c260)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_0                                                       (32'h260)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_1                                                   (32'h1001c264)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_1                                                       (32'h264)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_2                                                   (32'h1001c268)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_2                                                       (32'h268)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_3                                                   (32'h1001c26c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_3                                                       (32'h26c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_4                                                   (32'h1001c270)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_4                                                       (32'h270)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_5                                                   (32'h1001c274)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_5                                                       (32'h274)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_6                                                   (32'h1001c278)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_6                                                       (32'h278)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_7                                                   (32'h1001c27c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_7                                                       (32'h27c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_8                                                   (32'h1001c280)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_8                                                       (32'h280)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_9                                                   (32'h1001c284)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_9                                                       (32'h284)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_10                                                  (32'h1001c288)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_10                                                      (32'h288)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_11                                                  (32'h1001c28c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_1_11                                                      (32'h28c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_0                                                   (32'h1001c290)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_0                                                       (32'h290)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_1                                                   (32'h1001c294)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_1                                                       (32'h294)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_2                                                   (32'h1001c298)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_2                                                       (32'h298)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_3                                                   (32'h1001c29c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_3                                                       (32'h29c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_4                                                   (32'h1001c2a0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_4                                                       (32'h2a0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_5                                                   (32'h1001c2a4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_5                                                       (32'h2a4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_6                                                   (32'h1001c2a8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_6                                                       (32'h2a8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_7                                                   (32'h1001c2ac)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_7                                                       (32'h2ac)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_8                                                   (32'h1001c2b0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_8                                                       (32'h2b0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_9                                                   (32'h1001c2b4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_9                                                       (32'h2b4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_10                                                  (32'h1001c2b8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_10                                                      (32'h2b8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_11                                                  (32'h1001c2bc)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_2_11                                                      (32'h2bc)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_0                                                   (32'h1001c2c0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_0                                                       (32'h2c0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_1                                                   (32'h1001c2c4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_1                                                       (32'h2c4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_2                                                   (32'h1001c2c8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_2                                                       (32'h2c8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_3                                                   (32'h1001c2cc)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_3                                                       (32'h2cc)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_4                                                   (32'h1001c2d0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_4                                                       (32'h2d0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_5                                                   (32'h1001c2d4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_5                                                       (32'h2d4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_6                                                   (32'h1001c2d8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_6                                                       (32'h2d8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_7                                                   (32'h1001c2dc)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_7                                                       (32'h2dc)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_8                                                   (32'h1001c2e0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_8                                                       (32'h2e0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_9                                                   (32'h1001c2e4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_9                                                       (32'h2e4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_10                                                  (32'h1001c2e8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_10                                                      (32'h2e8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_11                                                  (32'h1001c2ec)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_3_11                                                      (32'h2ec)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_0                                                   (32'h1001c2f0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_0                                                       (32'h2f0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_1                                                   (32'h1001c2f4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_1                                                       (32'h2f4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_2                                                   (32'h1001c2f8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_2                                                       (32'h2f8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_3                                                   (32'h1001c2fc)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_3                                                       (32'h2fc)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_4                                                   (32'h1001c300)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_4                                                       (32'h300)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_5                                                   (32'h1001c304)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_5                                                       (32'h304)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_6                                                   (32'h1001c308)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_6                                                       (32'h308)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_7                                                   (32'h1001c30c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_7                                                       (32'h30c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_8                                                   (32'h1001c310)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_8                                                       (32'h310)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_9                                                   (32'h1001c314)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_9                                                       (32'h314)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_10                                                  (32'h1001c318)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_10                                                      (32'h318)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_11                                                  (32'h1001c31c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_4_11                                                      (32'h31c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_0                                                   (32'h1001c320)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_0                                                       (32'h320)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_1                                                   (32'h1001c324)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_1                                                       (32'h324)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_2                                                   (32'h1001c328)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_2                                                       (32'h328)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_3                                                   (32'h1001c32c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_3                                                       (32'h32c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_4                                                   (32'h1001c330)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_4                                                       (32'h330)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_5                                                   (32'h1001c334)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_5                                                       (32'h334)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_6                                                   (32'h1001c338)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_6                                                       (32'h338)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_7                                                   (32'h1001c33c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_7                                                       (32'h33c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_8                                                   (32'h1001c340)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_8                                                       (32'h340)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_9                                                   (32'h1001c344)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_9                                                       (32'h344)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_10                                                  (32'h1001c348)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_10                                                      (32'h348)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_11                                                  (32'h1001c34c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_5_11                                                      (32'h34c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_0                                                   (32'h1001c350)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_0                                                       (32'h350)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_1                                                   (32'h1001c354)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_1                                                       (32'h354)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_2                                                   (32'h1001c358)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_2                                                       (32'h358)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_3                                                   (32'h1001c35c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_3                                                       (32'h35c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_4                                                   (32'h1001c360)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_4                                                       (32'h360)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_5                                                   (32'h1001c364)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_5                                                       (32'h364)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_6                                                   (32'h1001c368)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_6                                                       (32'h368)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_7                                                   (32'h1001c36c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_7                                                       (32'h36c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_8                                                   (32'h1001c370)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_8                                                       (32'h370)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_9                                                   (32'h1001c374)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_9                                                       (32'h374)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_10                                                  (32'h1001c378)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_10                                                      (32'h378)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_11                                                  (32'h1001c37c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_6_11                                                      (32'h37c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_0                                                   (32'h1001c380)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_0                                                       (32'h380)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_1                                                   (32'h1001c384)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_1                                                       (32'h384)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_2                                                   (32'h1001c388)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_2                                                       (32'h388)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_3                                                   (32'h1001c38c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_3                                                       (32'h38c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_4                                                   (32'h1001c390)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_4                                                       (32'h390)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_5                                                   (32'h1001c394)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_5                                                       (32'h394)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_6                                                   (32'h1001c398)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_6                                                       (32'h398)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_7                                                   (32'h1001c39c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_7                                                       (32'h39c)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_8                                                   (32'h1001c3a0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_8                                                       (32'h3a0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_9                                                   (32'h1001c3a4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_9                                                       (32'h3a4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_10                                                  (32'h1001c3a8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_10                                                      (32'h3a8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_11                                                  (32'h1001c3ac)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_7_11                                                      (32'h3ac)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_0                                                   (32'h1001c3b0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_0                                                       (32'h3b0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_1                                                   (32'h1001c3b4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_1                                                       (32'h3b4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_2                                                   (32'h1001c3b8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_2                                                       (32'h3b8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_3                                                   (32'h1001c3bc)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_3                                                       (32'h3bc)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_4                                                   (32'h1001c3c0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_4                                                       (32'h3c0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_5                                                   (32'h1001c3c4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_5                                                       (32'h3c4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_6                                                   (32'h1001c3c8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_6                                                       (32'h3c8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_7                                                   (32'h1001c3cc)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_7                                                       (32'h3cc)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_8                                                   (32'h1001c3d0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_8                                                       (32'h3d0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_9                                                   (32'h1001c3d4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_9                                                       (32'h3d4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_10                                                  (32'h1001c3d8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_10                                                      (32'h3d8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_11                                                  (32'h1001c3dc)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_8_11                                                      (32'h3dc)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_0                                                   (32'h1001c3e0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_0                                                       (32'h3e0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_1                                                   (32'h1001c3e4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_1                                                       (32'h3e4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_2                                                   (32'h1001c3e8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_2                                                       (32'h3e8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_3                                                   (32'h1001c3ec)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_3                                                       (32'h3ec)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_4                                                   (32'h1001c3f0)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_4                                                       (32'h3f0)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_5                                                   (32'h1001c3f4)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_5                                                       (32'h3f4)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_6                                                   (32'h1001c3f8)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_6                                                       (32'h3f8)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_7                                                   (32'h1001c3fc)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_7                                                       (32'h3fc)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_8                                                   (32'h1001c400)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_8                                                       (32'h400)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_9                                                   (32'h1001c404)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_9                                                       (32'h404)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_10                                                  (32'h1001c408)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_10                                                      (32'h408)
`define CLP_DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_11                                                  (32'h1001c40c)
`define DV_REG_NONSTICKY_DATA_VAULT_ENTRY_9_11                                                      (32'h40c)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_0                                                (32'h1001c410)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_0                                                    (32'h410)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_0_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_0_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_1                                                (32'h1001c414)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_1                                                    (32'h414)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_1_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_1_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_2                                                (32'h1001c418)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_2                                                    (32'h418)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_2_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_2_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_3                                                (32'h1001c41c)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_3                                                    (32'h41c)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_3_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_3_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_4                                                (32'h1001c420)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_4                                                    (32'h420)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_4_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_4_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_5                                                (32'h1001c424)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_5                                                    (32'h424)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_5_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_5_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_6                                                (32'h1001c428)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_6                                                    (32'h428)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_6_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_6_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_7                                                (32'h1001c42c)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_7                                                    (32'h42c)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_7_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_7_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_8                                                (32'h1001c430)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_8                                                    (32'h430)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_8_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_8_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_9                                                (32'h1001c434)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_9                                                    (32'h434)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_9_LOCK_ENTRY_LOW                                     (0)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREGCTRL_9_LOCK_ENTRY_MASK                                    (32'h1)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_0                                                    (32'h1001c438)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_0                                                        (32'h438)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_1                                                    (32'h1001c43c)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_1                                                        (32'h43c)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_2                                                    (32'h1001c440)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_2                                                        (32'h440)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_3                                                    (32'h1001c444)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_3                                                        (32'h444)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_4                                                    (32'h1001c448)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_4                                                        (32'h448)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_5                                                    (32'h1001c44c)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_5                                                        (32'h44c)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_6                                                    (32'h1001c450)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_6                                                        (32'h450)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_7                                                    (32'h1001c454)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_7                                                        (32'h454)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_8                                                    (32'h1001c458)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_8                                                        (32'h458)
`define CLP_DV_REG_NONSTICKYLOCKABLESCRATCHREG_9                                                    (32'h1001c45c)
`define DV_REG_NONSTICKYLOCKABLESCRATCHREG_9                                                        (32'h45c)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_0                                                     (32'h1001c460)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_0                                                         (32'h460)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_1                                                     (32'h1001c464)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_1                                                         (32'h464)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_2                                                     (32'h1001c468)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_2                                                         (32'h468)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_3                                                     (32'h1001c46c)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_3                                                         (32'h46c)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_4                                                     (32'h1001c470)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_4                                                         (32'h470)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_5                                                     (32'h1001c474)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_5                                                         (32'h474)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_6                                                     (32'h1001c478)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_6                                                         (32'h478)
`define CLP_DV_REG_NONSTICKYGENERICSCRATCHREG_7                                                     (32'h1001c47c)
`define DV_REG_NONSTICKYGENERICSCRATCHREG_7                                                         (32'h47c)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0                                                   (32'h1001c480)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0                                                       (32'h480)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_0_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1                                                   (32'h1001c484)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1                                                       (32'h484)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_1_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2                                                   (32'h1001c488)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2                                                       (32'h488)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_2_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3                                                   (32'h1001c48c)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3                                                       (32'h48c)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_3_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4                                                   (32'h1001c490)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4                                                       (32'h490)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_4_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5                                                   (32'h1001c494)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5                                                       (32'h494)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_5_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6                                                   (32'h1001c498)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6                                                       (32'h498)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_6_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7                                                   (32'h1001c49c)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7                                                       (32'h49c)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7_LOCK_ENTRY_LOW                                        (0)
`define DV_REG_STICKYLOCKABLESCRATCHREGCTRL_7_LOCK_ENTRY_MASK                                       (32'h1)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_0                                                       (32'h1001c4a0)
`define DV_REG_STICKYLOCKABLESCRATCHREG_0                                                           (32'h4a0)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_1                                                       (32'h1001c4a4)
`define DV_REG_STICKYLOCKABLESCRATCHREG_1                                                           (32'h4a4)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_2                                                       (32'h1001c4a8)
`define DV_REG_STICKYLOCKABLESCRATCHREG_2                                                           (32'h4a8)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_3                                                       (32'h1001c4ac)
`define DV_REG_STICKYLOCKABLESCRATCHREG_3                                                           (32'h4ac)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_4                                                       (32'h1001c4b0)
`define DV_REG_STICKYLOCKABLESCRATCHREG_4                                                           (32'h4b0)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_5                                                       (32'h1001c4b4)
`define DV_REG_STICKYLOCKABLESCRATCHREG_5                                                           (32'h4b4)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_6                                                       (32'h1001c4b8)
`define DV_REG_STICKYLOCKABLESCRATCHREG_6                                                           (32'h4b8)
`define CLP_DV_REG_STICKYLOCKABLESCRATCHREG_7                                                       (32'h1001c4bc)
`define DV_REG_STICKYLOCKABLESCRATCHREG_7                                                           (32'h4bc)
`define CLP_SHA512_REG_BASE_ADDR                                                                    (32'h10020000)
`define CLP_SHA512_REG_SHA512_NAME_0                                                                (32'h10020000)
`define SHA512_REG_SHA512_NAME_0                                                                    (32'h0)
`define CLP_SHA512_REG_SHA512_NAME_1                                                                (32'h10020004)
`define SHA512_REG_SHA512_NAME_1                                                                    (32'h4)
`define CLP_SHA512_REG_SHA512_VERSION_0                                                             (32'h10020008)
`define SHA512_REG_SHA512_VERSION_0                                                                 (32'h8)
`define CLP_SHA512_REG_SHA512_VERSION_1                                                             (32'h1002000c)
`define SHA512_REG_SHA512_VERSION_1                                                                 (32'hc)
`define CLP_SHA512_REG_SHA512_CTRL                                                                  (32'h10020010)
`define SHA512_REG_SHA512_CTRL                                                                      (32'h10)
`define SHA512_REG_SHA512_CTRL_INIT_LOW                                                             (0)
`define SHA512_REG_SHA512_CTRL_INIT_MASK                                                            (32'h1)
`define SHA512_REG_SHA512_CTRL_NEXT_LOW                                                             (1)
`define SHA512_REG_SHA512_CTRL_NEXT_MASK                                                            (32'h2)
`define SHA512_REG_SHA512_CTRL_MODE_LOW                                                             (2)
`define SHA512_REG_SHA512_CTRL_MODE_MASK                                                            (32'hc)
`define SHA512_REG_SHA512_CTRL_ZEROIZE_LOW                                                          (4)
`define SHA512_REG_SHA512_CTRL_ZEROIZE_MASK                                                         (32'h10)
`define SHA512_REG_SHA512_CTRL_LAST_LOW                                                             (5)
`define SHA512_REG_SHA512_CTRL_LAST_MASK                                                            (32'h20)
`define CLP_SHA512_REG_SHA512_STATUS                                                                (32'h10020018)
`define SHA512_REG_SHA512_STATUS                                                                    (32'h18)
`define SHA512_REG_SHA512_STATUS_READY_LOW                                                          (0)
`define SHA512_REG_SHA512_STATUS_READY_MASK                                                         (32'h1)
`define SHA512_REG_SHA512_STATUS_VALID_LOW                                                          (1)
`define SHA512_REG_SHA512_STATUS_VALID_MASK                                                         (32'h2)
`define CLP_SHA512_REG_SHA512_BLOCK_0                                                               (32'h10020080)
`define SHA512_REG_SHA512_BLOCK_0                                                                   (32'h80)
`define CLP_SHA512_REG_SHA512_BLOCK_1                                                               (32'h10020084)
`define SHA512_REG_SHA512_BLOCK_1                                                                   (32'h84)
`define CLP_SHA512_REG_SHA512_BLOCK_2                                                               (32'h10020088)
`define SHA512_REG_SHA512_BLOCK_2                                                                   (32'h88)
`define CLP_SHA512_REG_SHA512_BLOCK_3                                                               (32'h1002008c)
`define SHA512_REG_SHA512_BLOCK_3                                                                   (32'h8c)
`define CLP_SHA512_REG_SHA512_BLOCK_4                                                               (32'h10020090)
`define SHA512_REG_SHA512_BLOCK_4                                                                   (32'h90)
`define CLP_SHA512_REG_SHA512_BLOCK_5                                                               (32'h10020094)
`define SHA512_REG_SHA512_BLOCK_5                                                                   (32'h94)
`define CLP_SHA512_REG_SHA512_BLOCK_6                                                               (32'h10020098)
`define SHA512_REG_SHA512_BLOCK_6                                                                   (32'h98)
`define CLP_SHA512_REG_SHA512_BLOCK_7                                                               (32'h1002009c)
`define SHA512_REG_SHA512_BLOCK_7                                                                   (32'h9c)
`define CLP_SHA512_REG_SHA512_BLOCK_8                                                               (32'h100200a0)
`define SHA512_REG_SHA512_BLOCK_8                                                                   (32'ha0)
`define CLP_SHA512_REG_SHA512_BLOCK_9                                                               (32'h100200a4)
`define SHA512_REG_SHA512_BLOCK_9                                                                   (32'ha4)
`define CLP_SHA512_REG_SHA512_BLOCK_10                                                              (32'h100200a8)
`define SHA512_REG_SHA512_BLOCK_10                                                                  (32'ha8)
`define CLP_SHA512_REG_SHA512_BLOCK_11                                                              (32'h100200ac)
`define SHA512_REG_SHA512_BLOCK_11                                                                  (32'hac)
`define CLP_SHA512_REG_SHA512_BLOCK_12                                                              (32'h100200b0)
`define SHA512_REG_SHA512_BLOCK_12                                                                  (32'hb0)
`define CLP_SHA512_REG_SHA512_BLOCK_13                                                              (32'h100200b4)
`define SHA512_REG_SHA512_BLOCK_13                                                                  (32'hb4)
`define CLP_SHA512_REG_SHA512_BLOCK_14                                                              (32'h100200b8)
`define SHA512_REG_SHA512_BLOCK_14                                                                  (32'hb8)
`define CLP_SHA512_REG_SHA512_BLOCK_15                                                              (32'h100200bc)
`define SHA512_REG_SHA512_BLOCK_15                                                                  (32'hbc)
`define CLP_SHA512_REG_SHA512_BLOCK_16                                                              (32'h100200c0)
`define SHA512_REG_SHA512_BLOCK_16                                                                  (32'hc0)
`define CLP_SHA512_REG_SHA512_BLOCK_17                                                              (32'h100200c4)
`define SHA512_REG_SHA512_BLOCK_17                                                                  (32'hc4)
`define CLP_SHA512_REG_SHA512_BLOCK_18                                                              (32'h100200c8)
`define SHA512_REG_SHA512_BLOCK_18                                                                  (32'hc8)
`define CLP_SHA512_REG_SHA512_BLOCK_19                                                              (32'h100200cc)
`define SHA512_REG_SHA512_BLOCK_19                                                                  (32'hcc)
`define CLP_SHA512_REG_SHA512_BLOCK_20                                                              (32'h100200d0)
`define SHA512_REG_SHA512_BLOCK_20                                                                  (32'hd0)
`define CLP_SHA512_REG_SHA512_BLOCK_21                                                              (32'h100200d4)
`define SHA512_REG_SHA512_BLOCK_21                                                                  (32'hd4)
`define CLP_SHA512_REG_SHA512_BLOCK_22                                                              (32'h100200d8)
`define SHA512_REG_SHA512_BLOCK_22                                                                  (32'hd8)
`define CLP_SHA512_REG_SHA512_BLOCK_23                                                              (32'h100200dc)
`define SHA512_REG_SHA512_BLOCK_23                                                                  (32'hdc)
`define CLP_SHA512_REG_SHA512_BLOCK_24                                                              (32'h100200e0)
`define SHA512_REG_SHA512_BLOCK_24                                                                  (32'he0)
`define CLP_SHA512_REG_SHA512_BLOCK_25                                                              (32'h100200e4)
`define SHA512_REG_SHA512_BLOCK_25                                                                  (32'he4)
`define CLP_SHA512_REG_SHA512_BLOCK_26                                                              (32'h100200e8)
`define SHA512_REG_SHA512_BLOCK_26                                                                  (32'he8)
`define CLP_SHA512_REG_SHA512_BLOCK_27                                                              (32'h100200ec)
`define SHA512_REG_SHA512_BLOCK_27                                                                  (32'hec)
`define CLP_SHA512_REG_SHA512_BLOCK_28                                                              (32'h100200f0)
`define SHA512_REG_SHA512_BLOCK_28                                                                  (32'hf0)
`define CLP_SHA512_REG_SHA512_BLOCK_29                                                              (32'h100200f4)
`define SHA512_REG_SHA512_BLOCK_29                                                                  (32'hf4)
`define CLP_SHA512_REG_SHA512_BLOCK_30                                                              (32'h100200f8)
`define SHA512_REG_SHA512_BLOCK_30                                                                  (32'hf8)
`define CLP_SHA512_REG_SHA512_BLOCK_31                                                              (32'h100200fc)
`define SHA512_REG_SHA512_BLOCK_31                                                                  (32'hfc)
`define CLP_SHA512_REG_SHA512_DIGEST_0                                                              (32'h10020100)
`define SHA512_REG_SHA512_DIGEST_0                                                                  (32'h100)
`define CLP_SHA512_REG_SHA512_DIGEST_1                                                              (32'h10020104)
`define SHA512_REG_SHA512_DIGEST_1                                                                  (32'h104)
`define CLP_SHA512_REG_SHA512_DIGEST_2                                                              (32'h10020108)
`define SHA512_REG_SHA512_DIGEST_2                                                                  (32'h108)
`define CLP_SHA512_REG_SHA512_DIGEST_3                                                              (32'h1002010c)
`define SHA512_REG_SHA512_DIGEST_3                                                                  (32'h10c)
`define CLP_SHA512_REG_SHA512_DIGEST_4                                                              (32'h10020110)
`define SHA512_REG_SHA512_DIGEST_4                                                                  (32'h110)
`define CLP_SHA512_REG_SHA512_DIGEST_5                                                              (32'h10020114)
`define SHA512_REG_SHA512_DIGEST_5                                                                  (32'h114)
`define CLP_SHA512_REG_SHA512_DIGEST_6                                                              (32'h10020118)
`define SHA512_REG_SHA512_DIGEST_6                                                                  (32'h118)
`define CLP_SHA512_REG_SHA512_DIGEST_7                                                              (32'h1002011c)
`define SHA512_REG_SHA512_DIGEST_7                                                                  (32'h11c)
`define CLP_SHA512_REG_SHA512_DIGEST_8                                                              (32'h10020120)
`define SHA512_REG_SHA512_DIGEST_8                                                                  (32'h120)
`define CLP_SHA512_REG_SHA512_DIGEST_9                                                              (32'h10020124)
`define SHA512_REG_SHA512_DIGEST_9                                                                  (32'h124)
`define CLP_SHA512_REG_SHA512_DIGEST_10                                                             (32'h10020128)
`define SHA512_REG_SHA512_DIGEST_10                                                                 (32'h128)
`define CLP_SHA512_REG_SHA512_DIGEST_11                                                             (32'h1002012c)
`define SHA512_REG_SHA512_DIGEST_11                                                                 (32'h12c)
`define CLP_SHA512_REG_SHA512_DIGEST_12                                                             (32'h10020130)
`define SHA512_REG_SHA512_DIGEST_12                                                                 (32'h130)
`define CLP_SHA512_REG_SHA512_DIGEST_13                                                             (32'h10020134)
`define SHA512_REG_SHA512_DIGEST_13                                                                 (32'h134)
`define CLP_SHA512_REG_SHA512_DIGEST_14                                                             (32'h10020138)
`define SHA512_REG_SHA512_DIGEST_14                                                                 (32'h138)
`define CLP_SHA512_REG_SHA512_DIGEST_15                                                             (32'h1002013c)
`define SHA512_REG_SHA512_DIGEST_15                                                                 (32'h13c)
`define CLP_SHA512_REG_SHA512_VAULT_RD_CTRL                                                         (32'h10020600)
`define SHA512_REG_SHA512_VAULT_RD_CTRL                                                             (32'h600)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_READ_EN_LOW                                                 (0)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_READ_EN_MASK                                                (32'h1)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_READ_ENTRY_LOW                                              (1)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_READ_ENTRY_MASK                                             (32'h3e)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_PCR_HASH_EXTEND_LOW                                         (6)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_PCR_HASH_EXTEND_MASK                                        (32'h40)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_RSVD_LOW                                                    (7)
`define SHA512_REG_SHA512_VAULT_RD_CTRL_RSVD_MASK                                                   (32'hffffff80)
`define CLP_SHA512_REG_SHA512_VAULT_RD_STATUS                                                       (32'h10020604)
`define SHA512_REG_SHA512_VAULT_RD_STATUS                                                           (32'h604)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_READY_LOW                                                 (0)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_READY_MASK                                                (32'h1)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_VALID_LOW                                                 (1)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_VALID_MASK                                                (32'h2)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_ERROR_LOW                                                 (2)
`define SHA512_REG_SHA512_VAULT_RD_STATUS_ERROR_MASK                                                (32'h3fc)
`define CLP_SHA512_REG_SHA512_KV_WR_CTRL                                                            (32'h10020608)
`define SHA512_REG_SHA512_KV_WR_CTRL                                                                (32'h608)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_EN_LOW                                                   (0)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_EN_MASK                                                  (32'h1)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_ENTRY_LOW                                                (1)
`define SHA512_REG_SHA512_KV_WR_CTRL_WRITE_ENTRY_MASK                                               (32'h3e)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_KEY_DEST_VALID_LOW                                        (6)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_KEY_DEST_VALID_MASK                                       (32'h40)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_LOW                                      (7)
`define SHA512_REG_SHA512_KV_WR_CTRL_HMAC_BLOCK_DEST_VALID_MASK                                     (32'h80)
`define SHA512_REG_SHA512_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_LOW                                       (8)
`define SHA512_REG_SHA512_KV_WR_CTRL_SHA_BLOCK_DEST_VALID_MASK                                      (32'h100)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_PKEY_DEST_VALID_LOW                                        (9)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_PKEY_DEST_VALID_MASK                                       (32'h200)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_SEED_DEST_VALID_LOW                                        (10)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_SEED_DEST_VALID_MASK                                       (32'h400)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_MSG_DEST_VALID_LOW                                         (11)
`define SHA512_REG_SHA512_KV_WR_CTRL_ECC_MSG_DEST_VALID_MASK                                        (32'h800)
`define SHA512_REG_SHA512_KV_WR_CTRL_RSVD_LOW                                                       (12)
`define SHA512_REG_SHA512_KV_WR_CTRL_RSVD_MASK                                                      (32'hfffff000)
`define CLP_SHA512_REG_SHA512_KV_WR_STATUS                                                          (32'h1002060c)
`define SHA512_REG_SHA512_KV_WR_STATUS                                                              (32'h60c)
`define SHA512_REG_SHA512_KV_WR_STATUS_READY_LOW                                                    (0)
`define SHA512_REG_SHA512_KV_WR_STATUS_READY_MASK                                                   (32'h1)
`define SHA512_REG_SHA512_KV_WR_STATUS_VALID_LOW                                                    (1)
`define SHA512_REG_SHA512_KV_WR_STATUS_VALID_MASK                                                   (32'h2)
`define SHA512_REG_SHA512_KV_WR_STATUS_ERROR_LOW                                                    (2)
`define SHA512_REG_SHA512_KV_WR_STATUS_ERROR_MASK                                                   (32'h3fc)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_NONCE                                                    (32'h10020610)
`define SHA512_REG_SHA512_GEN_PCR_HASH_NONCE                                                        (32'h610)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_CTRL                                                     (32'h10020614)
`define SHA512_REG_SHA512_GEN_PCR_HASH_CTRL                                                         (32'h614)
`define SHA512_REG_SHA512_GEN_PCR_HASH_CTRL_START_LOW                                               (0)
`define SHA512_REG_SHA512_GEN_PCR_HASH_CTRL_START_MASK                                              (32'h1)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_STATUS                                                   (32'h10020618)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS                                                       (32'h618)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS_READY_LOW                                             (0)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS_READY_MASK                                            (32'h1)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS_VALID_LOW                                             (1)
`define SHA512_REG_SHA512_GEN_PCR_HASH_STATUS_VALID_MASK                                            (32'h2)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_0                                                 (32'h1002061c)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_0                                                     (32'h61c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_1                                                 (32'h10020620)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_1                                                     (32'h620)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_2                                                 (32'h10020624)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_2                                                     (32'h624)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_3                                                 (32'h10020628)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_3                                                     (32'h628)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_4                                                 (32'h1002062c)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_4                                                     (32'h62c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_5                                                 (32'h10020630)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_5                                                     (32'h630)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_6                                                 (32'h10020634)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_6                                                     (32'h634)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_7                                                 (32'h10020638)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_7                                                     (32'h638)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_8                                                 (32'h1002063c)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_8                                                     (32'h63c)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_9                                                 (32'h10020640)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_9                                                     (32'h640)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_10                                                (32'h10020644)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_10                                                    (32'h644)
`define CLP_SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_11                                                (32'h10020648)
`define SHA512_REG_SHA512_GEN_PCR_HASH_DIGEST_11                                                    (32'h648)
`define CLP_SHA512_REG_INTR_BLOCK_RF_START                                                          (32'h10020800)
`define CLP_SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h10020800)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                   (32'h800)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                      (0)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                     (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                      (1)
`define SHA512_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                     (32'h2)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h10020804)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                    (32'h804)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                      (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                     (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                      (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                     (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                      (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                     (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                      (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                     (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h10020808)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                    (32'h808)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                              (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                             (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h1002080c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                (32'h80c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h10020810)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                (32'h810)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h10020814)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                              (32'h814)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                               (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                              (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                               (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                              (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                               (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                              (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                               (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                              (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h10020818)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                              (32'h818)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                       (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                      (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h1002081c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                  (32'h81c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                  (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                 (32'h1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                  (1)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                 (32'h2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                  (2)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                 (32'h4)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                  (3)
`define SHA512_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                 (32'h8)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h10020820)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                  (32'h820)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                          (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                         (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h10020900)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                (32'h900)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h10020904)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                (32'h904)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h10020908)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                (32'h908)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h1002090c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                (32'h90c)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h10020980)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                        (32'h980)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'h10020a00)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                           (32'ha00)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'h10020a04)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                           (32'ha04)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'h10020a08)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                           (32'ha08)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'h10020a0c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                           (32'ha0c)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA512_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'h10020a10)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                   (32'ha10)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SHA512_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_SHA256_REG_BASE_ADDR                                                                    (32'h10028000)
`define CLP_SHA256_REG_SHA256_NAME_0                                                                (32'h10028000)
`define SHA256_REG_SHA256_NAME_0                                                                    (32'h0)
`define CLP_SHA256_REG_SHA256_NAME_1                                                                (32'h10028004)
`define SHA256_REG_SHA256_NAME_1                                                                    (32'h4)
`define CLP_SHA256_REG_SHA256_VERSION_0                                                             (32'h10028008)
`define SHA256_REG_SHA256_VERSION_0                                                                 (32'h8)
`define CLP_SHA256_REG_SHA256_VERSION_1                                                             (32'h1002800c)
`define SHA256_REG_SHA256_VERSION_1                                                                 (32'hc)
`define CLP_SHA256_REG_SHA256_CTRL                                                                  (32'h10028010)
`define SHA256_REG_SHA256_CTRL                                                                      (32'h10)
`define SHA256_REG_SHA256_CTRL_INIT_LOW                                                             (0)
`define SHA256_REG_SHA256_CTRL_INIT_MASK                                                            (32'h1)
`define SHA256_REG_SHA256_CTRL_NEXT_LOW                                                             (1)
`define SHA256_REG_SHA256_CTRL_NEXT_MASK                                                            (32'h2)
`define SHA256_REG_SHA256_CTRL_MODE_LOW                                                             (2)
`define SHA256_REG_SHA256_CTRL_MODE_MASK                                                            (32'h4)
`define SHA256_REG_SHA256_CTRL_ZEROIZE_LOW                                                          (3)
`define SHA256_REG_SHA256_CTRL_ZEROIZE_MASK                                                         (32'h8)
`define CLP_SHA256_REG_SHA256_STATUS                                                                (32'h10028018)
`define SHA256_REG_SHA256_STATUS                                                                    (32'h18)
`define SHA256_REG_SHA256_STATUS_READY_LOW                                                          (0)
`define SHA256_REG_SHA256_STATUS_READY_MASK                                                         (32'h1)
`define SHA256_REG_SHA256_STATUS_VALID_LOW                                                          (1)
`define SHA256_REG_SHA256_STATUS_VALID_MASK                                                         (32'h2)
`define CLP_SHA256_REG_SHA256_BLOCK_0                                                               (32'h10028080)
`define SHA256_REG_SHA256_BLOCK_0                                                                   (32'h80)
`define CLP_SHA256_REG_SHA256_BLOCK_1                                                               (32'h10028084)
`define SHA256_REG_SHA256_BLOCK_1                                                                   (32'h84)
`define CLP_SHA256_REG_SHA256_BLOCK_2                                                               (32'h10028088)
`define SHA256_REG_SHA256_BLOCK_2                                                                   (32'h88)
`define CLP_SHA256_REG_SHA256_BLOCK_3                                                               (32'h1002808c)
`define SHA256_REG_SHA256_BLOCK_3                                                                   (32'h8c)
`define CLP_SHA256_REG_SHA256_BLOCK_4                                                               (32'h10028090)
`define SHA256_REG_SHA256_BLOCK_4                                                                   (32'h90)
`define CLP_SHA256_REG_SHA256_BLOCK_5                                                               (32'h10028094)
`define SHA256_REG_SHA256_BLOCK_5                                                                   (32'h94)
`define CLP_SHA256_REG_SHA256_BLOCK_6                                                               (32'h10028098)
`define SHA256_REG_SHA256_BLOCK_6                                                                   (32'h98)
`define CLP_SHA256_REG_SHA256_BLOCK_7                                                               (32'h1002809c)
`define SHA256_REG_SHA256_BLOCK_7                                                                   (32'h9c)
`define CLP_SHA256_REG_SHA256_BLOCK_8                                                               (32'h100280a0)
`define SHA256_REG_SHA256_BLOCK_8                                                                   (32'ha0)
`define CLP_SHA256_REG_SHA256_BLOCK_9                                                               (32'h100280a4)
`define SHA256_REG_SHA256_BLOCK_9                                                                   (32'ha4)
`define CLP_SHA256_REG_SHA256_BLOCK_10                                                              (32'h100280a8)
`define SHA256_REG_SHA256_BLOCK_10                                                                  (32'ha8)
`define CLP_SHA256_REG_SHA256_BLOCK_11                                                              (32'h100280ac)
`define SHA256_REG_SHA256_BLOCK_11                                                                  (32'hac)
`define CLP_SHA256_REG_SHA256_BLOCK_12                                                              (32'h100280b0)
`define SHA256_REG_SHA256_BLOCK_12                                                                  (32'hb0)
`define CLP_SHA256_REG_SHA256_BLOCK_13                                                              (32'h100280b4)
`define SHA256_REG_SHA256_BLOCK_13                                                                  (32'hb4)
`define CLP_SHA256_REG_SHA256_BLOCK_14                                                              (32'h100280b8)
`define SHA256_REG_SHA256_BLOCK_14                                                                  (32'hb8)
`define CLP_SHA256_REG_SHA256_BLOCK_15                                                              (32'h100280bc)
`define SHA256_REG_SHA256_BLOCK_15                                                                  (32'hbc)
`define CLP_SHA256_REG_SHA256_DIGEST_0                                                              (32'h10028100)
`define SHA256_REG_SHA256_DIGEST_0                                                                  (32'h100)
`define CLP_SHA256_REG_SHA256_DIGEST_1                                                              (32'h10028104)
`define SHA256_REG_SHA256_DIGEST_1                                                                  (32'h104)
`define CLP_SHA256_REG_SHA256_DIGEST_2                                                              (32'h10028108)
`define SHA256_REG_SHA256_DIGEST_2                                                                  (32'h108)
`define CLP_SHA256_REG_SHA256_DIGEST_3                                                              (32'h1002810c)
`define SHA256_REG_SHA256_DIGEST_3                                                                  (32'h10c)
`define CLP_SHA256_REG_SHA256_DIGEST_4                                                              (32'h10028110)
`define SHA256_REG_SHA256_DIGEST_4                                                                  (32'h110)
`define CLP_SHA256_REG_SHA256_DIGEST_5                                                              (32'h10028114)
`define SHA256_REG_SHA256_DIGEST_5                                                                  (32'h114)
`define CLP_SHA256_REG_SHA256_DIGEST_6                                                              (32'h10028118)
`define SHA256_REG_SHA256_DIGEST_6                                                                  (32'h118)
`define CLP_SHA256_REG_SHA256_DIGEST_7                                                              (32'h1002811c)
`define SHA256_REG_SHA256_DIGEST_7                                                                  (32'h11c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_START                                                          (32'h10028800)
`define CLP_SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h10028800)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                   (32'h800)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                      (0)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                     (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                      (1)
`define SHA256_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                     (32'h2)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h10028804)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                    (32'h804)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                      (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                     (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                      (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                     (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                      (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                     (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                      (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                     (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h10028808)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                    (32'h808)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                              (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                             (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h1002880c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                                (32'h80c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h10028810)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                                (32'h810)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                    (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                   (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h10028814)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                              (32'h814)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                               (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                              (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                               (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                              (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                               (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                              (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                               (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                              (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h10028818)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                              (32'h818)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                       (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                      (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h1002881c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                  (32'h81c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                                  (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                                 (32'h1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                                  (1)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                                 (32'h2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                                  (2)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                                 (32'h4)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                                  (3)
`define SHA256_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                                 (32'h8)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h10028820)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                  (32'h820)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                          (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                         (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h10028900)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                                (32'h900)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h10028904)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                                (32'h904)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h10028908)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                                (32'h908)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h1002890c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                                (32'h90c)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h10028980)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                        (32'h980)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'h10028a00)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                           (32'ha00)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'h10028a04)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                           (32'ha04)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'h10028a08)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                           (32'ha08)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'h10028a0c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                           (32'ha0c)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                                 (0)
`define SHA256_REG_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                                (32'h1)
`define CLP_SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'h10028a10)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                                   (32'ha10)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SHA256_REG_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_MBOX_CSR_BASE_ADDR                                                                      (32'h30020000)
`define CLP_MBOX_CSR_MBOX_LOCK                                                                      (32'h30020000)
`define MBOX_CSR_MBOX_LOCK                                                                          (32'h0)
`define MBOX_CSR_MBOX_LOCK_LOCK_LOW                                                                 (0)
`define MBOX_CSR_MBOX_LOCK_LOCK_MASK                                                                (32'h1)
`define CLP_MBOX_CSR_MBOX_USER                                                                      (32'h30020004)
`define MBOX_CSR_MBOX_USER                                                                          (32'h4)
`define CLP_MBOX_CSR_MBOX_CMD                                                                       (32'h30020008)
`define MBOX_CSR_MBOX_CMD                                                                           (32'h8)
`define CLP_MBOX_CSR_MBOX_DLEN                                                                      (32'h3002000c)
`define MBOX_CSR_MBOX_DLEN                                                                          (32'hc)
`define CLP_MBOX_CSR_MBOX_DATAIN                                                                    (32'h30020010)
`define MBOX_CSR_MBOX_DATAIN                                                                        (32'h10)
`define CLP_MBOX_CSR_MBOX_DATAOUT                                                                   (32'h30020014)
`define MBOX_CSR_MBOX_DATAOUT                                                                       (32'h14)
`define CLP_MBOX_CSR_MBOX_EXECUTE                                                                   (32'h30020018)
`define MBOX_CSR_MBOX_EXECUTE                                                                       (32'h18)
`define MBOX_CSR_MBOX_EXECUTE_EXECUTE_LOW                                                           (0)
`define MBOX_CSR_MBOX_EXECUTE_EXECUTE_MASK                                                          (32'h1)
`define CLP_MBOX_CSR_MBOX_STATUS                                                                    (32'h3002001c)
`define MBOX_CSR_MBOX_STATUS                                                                        (32'h1c)
`define MBOX_CSR_MBOX_STATUS_STATUS_LOW                                                             (0)
`define MBOX_CSR_MBOX_STATUS_STATUS_MASK                                                            (32'hf)
`define MBOX_CSR_MBOX_STATUS_ECC_SINGLE_ERROR_LOW                                                   (4)
`define MBOX_CSR_MBOX_STATUS_ECC_SINGLE_ERROR_MASK                                                  (32'h10)
`define MBOX_CSR_MBOX_STATUS_ECC_DOUBLE_ERROR_LOW                                                   (5)
`define MBOX_CSR_MBOX_STATUS_ECC_DOUBLE_ERROR_MASK                                                  (32'h20)
`define MBOX_CSR_MBOX_STATUS_MBOX_FSM_PS_LOW                                                        (6)
`define MBOX_CSR_MBOX_STATUS_MBOX_FSM_PS_MASK                                                       (32'h1c0)
`define MBOX_CSR_MBOX_STATUS_SOC_HAS_LOCK_LOW                                                       (9)
`define MBOX_CSR_MBOX_STATUS_SOC_HAS_LOCK_MASK                                                      (32'h200)
`define CLP_MBOX_CSR_MBOX_UNLOCK                                                                    (32'h30020020)
`define MBOX_CSR_MBOX_UNLOCK                                                                        (32'h20)
`define MBOX_CSR_MBOX_UNLOCK_UNLOCK_LOW                                                             (0)
`define MBOX_CSR_MBOX_UNLOCK_UNLOCK_MASK                                                            (32'h1)
`define CLP_SHA512_ACC_CSR_BASE_ADDR                                                                (32'h30021000)
`define CLP_SHA512_ACC_CSR_LOCK                                                                     (32'h30021000)
`define SHA512_ACC_CSR_LOCK                                                                         (32'h0)
`define SHA512_ACC_CSR_LOCK_LOCK_LOW                                                                (0)
`define SHA512_ACC_CSR_LOCK_LOCK_MASK                                                               (32'h1)
`define CLP_SHA512_ACC_CSR_USER                                                                     (32'h30021004)
`define SHA512_ACC_CSR_USER                                                                         (32'h4)
`define CLP_SHA512_ACC_CSR_MODE                                                                     (32'h30021008)
`define SHA512_ACC_CSR_MODE                                                                         (32'h8)
`define SHA512_ACC_CSR_MODE_MODE_LOW                                                                (0)
`define SHA512_ACC_CSR_MODE_MODE_MASK                                                               (32'h3)
`define SHA512_ACC_CSR_MODE_ENDIAN_TOGGLE_LOW                                                       (2)
`define SHA512_ACC_CSR_MODE_ENDIAN_TOGGLE_MASK                                                      (32'h4)
`define CLP_SHA512_ACC_CSR_START_ADDRESS                                                            (32'h3002100c)
`define SHA512_ACC_CSR_START_ADDRESS                                                                (32'hc)
`define CLP_SHA512_ACC_CSR_DLEN                                                                     (32'h30021010)
`define SHA512_ACC_CSR_DLEN                                                                         (32'h10)
`define CLP_SHA512_ACC_CSR_DATAIN                                                                   (32'h30021014)
`define SHA512_ACC_CSR_DATAIN                                                                       (32'h14)
`define CLP_SHA512_ACC_CSR_EXECUTE                                                                  (32'h30021018)
`define SHA512_ACC_CSR_EXECUTE                                                                      (32'h18)
`define SHA512_ACC_CSR_EXECUTE_EXECUTE_LOW                                                          (0)
`define SHA512_ACC_CSR_EXECUTE_EXECUTE_MASK                                                         (32'h1)
`define CLP_SHA512_ACC_CSR_STATUS                                                                   (32'h3002101c)
`define SHA512_ACC_CSR_STATUS                                                                       (32'h1c)
`define SHA512_ACC_CSR_STATUS_VALID_LOW                                                             (0)
`define SHA512_ACC_CSR_STATUS_VALID_MASK                                                            (32'h1)
`define CLP_SHA512_ACC_CSR_DIGEST_0                                                                 (32'h30021020)
`define SHA512_ACC_CSR_DIGEST_0                                                                     (32'h20)
`define CLP_SHA512_ACC_CSR_DIGEST_1                                                                 (32'h30021024)
`define SHA512_ACC_CSR_DIGEST_1                                                                     (32'h24)
`define CLP_SHA512_ACC_CSR_DIGEST_2                                                                 (32'h30021028)
`define SHA512_ACC_CSR_DIGEST_2                                                                     (32'h28)
`define CLP_SHA512_ACC_CSR_DIGEST_3                                                                 (32'h3002102c)
`define SHA512_ACC_CSR_DIGEST_3                                                                     (32'h2c)
`define CLP_SHA512_ACC_CSR_DIGEST_4                                                                 (32'h30021030)
`define SHA512_ACC_CSR_DIGEST_4                                                                     (32'h30)
`define CLP_SHA512_ACC_CSR_DIGEST_5                                                                 (32'h30021034)
`define SHA512_ACC_CSR_DIGEST_5                                                                     (32'h34)
`define CLP_SHA512_ACC_CSR_DIGEST_6                                                                 (32'h30021038)
`define SHA512_ACC_CSR_DIGEST_6                                                                     (32'h38)
`define CLP_SHA512_ACC_CSR_DIGEST_7                                                                 (32'h3002103c)
`define SHA512_ACC_CSR_DIGEST_7                                                                     (32'h3c)
`define CLP_SHA512_ACC_CSR_DIGEST_8                                                                 (32'h30021040)
`define SHA512_ACC_CSR_DIGEST_8                                                                     (32'h40)
`define CLP_SHA512_ACC_CSR_DIGEST_9                                                                 (32'h30021044)
`define SHA512_ACC_CSR_DIGEST_9                                                                     (32'h44)
`define CLP_SHA512_ACC_CSR_DIGEST_10                                                                (32'h30021048)
`define SHA512_ACC_CSR_DIGEST_10                                                                    (32'h48)
`define CLP_SHA512_ACC_CSR_DIGEST_11                                                                (32'h3002104c)
`define SHA512_ACC_CSR_DIGEST_11                                                                    (32'h4c)
`define CLP_SHA512_ACC_CSR_DIGEST_12                                                                (32'h30021050)
`define SHA512_ACC_CSR_DIGEST_12                                                                    (32'h50)
`define CLP_SHA512_ACC_CSR_DIGEST_13                                                                (32'h30021054)
`define SHA512_ACC_CSR_DIGEST_13                                                                    (32'h54)
`define CLP_SHA512_ACC_CSR_DIGEST_14                                                                (32'h30021058)
`define SHA512_ACC_CSR_DIGEST_14                                                                    (32'h58)
`define CLP_SHA512_ACC_CSR_DIGEST_15                                                                (32'h3002105c)
`define SHA512_ACC_CSR_DIGEST_15                                                                    (32'h5c)
`define CLP_SHA512_ACC_CSR_CONTROL                                                                  (32'h30021060)
`define SHA512_ACC_CSR_CONTROL                                                                      (32'h60)
`define SHA512_ACC_CSR_CONTROL_ZEROIZE_LOW                                                          (0)
`define SHA512_ACC_CSR_CONTROL_ZEROIZE_MASK                                                         (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_START                                                      (32'h30021800)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                           (32'h30021800)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                               (32'h800)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                  (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                 (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                  (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                 (32'h2)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R                                            (32'h30021804)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                (32'h804)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_LOW                                  (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR0_EN_MASK                                 (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_LOW                                  (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR1_EN_MASK                                 (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_LOW                                  (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR2_EN_MASK                                 (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_LOW                                  (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR3_EN_MASK                                 (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                            (32'h30021808)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                (32'h808)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_LOW                          (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_DONE_EN_MASK                         (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                        (32'h3002180c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                            (32'h80c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                               (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                        (32'h30021810)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                            (32'h810)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                               (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                      (32'h30021814)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                          (32'h814)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_LOW                           (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR0_STS_MASK                          (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_LOW                           (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR1_STS_MASK                          (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_LOW                           (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR2_STS_MASK                          (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_LOW                           (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR3_STS_MASK                          (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                      (32'h30021818)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                          (32'h818)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_LOW                   (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_DONE_STS_MASK                  (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                          (32'h3002181c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                              (32'h81c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_LOW                              (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR0_TRIG_MASK                             (32'h1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_LOW                              (1)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR1_TRIG_MASK                             (32'h2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_LOW                              (2)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR2_TRIG_MASK                             (32'h4)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_LOW                              (3)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR3_TRIG_MASK                             (32'h8)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                          (32'h30021820)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                              (32'h820)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_LOW                      (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_DONE_TRIG_MASK                     (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                        (32'h30021900)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_R                                            (32'h900)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                        (32'h30021904)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_R                                            (32'h904)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                        (32'h30021908)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_R                                            (32'h908)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                        (32'h3002190c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_R                                            (32'h90c)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                (32'h30021980)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_R                                    (32'h980)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                   (32'h30021a00)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R                                       (32'ha00)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR0_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                   (32'h30021a04)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R                                       (32'ha04)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR1_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                   (32'h30021a08)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R                                       (32'ha08)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR2_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                   (32'h30021a0c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R                                       (32'ha0c)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_LOW                             (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_ERROR3_INTR_COUNT_INCR_R_PULSE_MASK                            (32'h1)
`define CLP_SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                           (32'h30021a10)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R                               (32'ha10)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_LOW                     (0)
`define SHA512_ACC_CSR_INTR_BLOCK_RF_NOTIF_CMD_DONE_INTR_COUNT_INCR_R_PULSE_MASK                    (32'h1)
`define CLP_SOC_IFC_REG_BASE_ADDR                                                                   (32'h30030000)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_FATAL                                                        (32'h30030000)
`define SOC_IFC_REG_CPTRA_HW_ERROR_FATAL                                                            (32'h0)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL                                                    (32'h30030004)
`define SOC_IFC_REG_CPTRA_HW_ERROR_NON_FATAL                                                        (32'h4)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_FATAL                                                        (32'h30030008)
`define SOC_IFC_REG_CPTRA_FW_ERROR_FATAL                                                            (32'h8)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_NON_FATAL                                                    (32'h3003000c)
`define SOC_IFC_REG_CPTRA_FW_ERROR_NON_FATAL                                                        (32'hc)
`define CLP_SOC_IFC_REG_CPTRA_HW_ERROR_ENC                                                          (32'h30030010)
`define SOC_IFC_REG_CPTRA_HW_ERROR_ENC                                                              (32'h10)
`define CLP_SOC_IFC_REG_CPTRA_FW_ERROR_ENC                                                          (32'h30030014)
`define SOC_IFC_REG_CPTRA_FW_ERROR_ENC                                                              (32'h14)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                              (32'h30030018)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_0                                                  (32'h18)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                              (32'h3003001c)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_1                                                  (32'h1c)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                              (32'h30030020)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_2                                                  (32'h20)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                              (32'h30030024)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_3                                                  (32'h24)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                              (32'h30030028)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_4                                                  (32'h28)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                              (32'h3003002c)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_5                                                  (32'h2c)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                              (32'h30030030)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_6                                                  (32'h30)
`define CLP_SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                              (32'h30030034)
`define SOC_IFC_REG_CPTRA_FW_EXTENDED_ERROR_INFO_7                                                  (32'h34)
`define CLP_SOC_IFC_REG_CPTRA_BOOT_STATUS                                                           (32'h30030038)
`define SOC_IFC_REG_CPTRA_BOOT_STATUS                                                               (32'h38)
`define CLP_SOC_IFC_REG_CPTRA_FLOW_STATUS                                                           (32'h3003003c)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS                                                               (32'h3c)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_STATUS_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_STATUS_MASK                                                   (32'hfffffff)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FW_LOW                                              (28)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FW_MASK                                             (32'h10000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_RUNTIME_LOW                                         (29)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_RUNTIME_MASK                                        (32'h20000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FUSES_LOW                                           (30)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_READY_FOR_FUSES_MASK                                          (32'h40000000)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_MAILBOX_FLOW_DONE_LOW                                         (31)
`define SOC_IFC_REG_CPTRA_FLOW_STATUS_MAILBOX_FLOW_DONE_MASK                                        (32'h80000000)
`define CLP_SOC_IFC_REG_CPTRA_RESET_REASON                                                          (32'h30030040)
`define SOC_IFC_REG_CPTRA_RESET_REASON                                                              (32'h40)
`define SOC_IFC_REG_CPTRA_RESET_REASON_FW_UPD_RESET_LOW                                             (0)
`define SOC_IFC_REG_CPTRA_RESET_REASON_FW_UPD_RESET_MASK                                            (32'h1)
`define SOC_IFC_REG_CPTRA_RESET_REASON_WARM_RESET_LOW                                               (1)
`define SOC_IFC_REG_CPTRA_RESET_REASON_WARM_RESET_MASK                                              (32'h2)
`define CLP_SOC_IFC_REG_CPTRA_SECURITY_STATE                                                        (32'h30030044)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE                                                            (32'h44)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEVICE_LIFECYCLE_LOW                                       (0)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEVICE_LIFECYCLE_MASK                                      (32'h3)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEBUG_LOCKED_LOW                                           (2)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_DEBUG_LOCKED_MASK                                          (32'h4)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_SCAN_MODE_LOW                                              (3)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_SCAN_MODE_MASK                                             (32'h8)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_RSVD_LOW                                                   (4)
`define SOC_IFC_REG_CPTRA_SECURITY_STATE_RSVD_MASK                                                  (32'hfffffff0)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_0                                                        (32'h30030048)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_0                                                            (32'h48)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_1                                                        (32'h3003004c)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_1                                                            (32'h4c)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_2                                                        (32'h30030050)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_2                                                            (32'h50)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_3                                                        (32'h30030054)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_3                                                            (32'h54)
`define CLP_SOC_IFC_REG_CPTRA_VALID_PAUSER_4                                                        (32'h30030058)
`define SOC_IFC_REG_CPTRA_VALID_PAUSER_4                                                            (32'h58)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_0                                                         (32'h3003005c)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_0                                                             (32'h5c)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_0_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_0_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_1                                                         (32'h30030060)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_1                                                             (32'h60)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_1_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_1_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_2                                                         (32'h30030064)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_2                                                             (32'h64)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_2_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_2_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_3                                                         (32'h30030068)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_3                                                             (32'h68)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_3_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_3_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_PAUSER_LOCK_4                                                         (32'h3003006c)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_4                                                             (32'h6c)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_4_LOCK_LOW                                                    (0)
`define SOC_IFC_REG_CPTRA_PAUSER_LOCK_4_LOCK_MASK                                                   (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_VALID_PAUSER                                                     (32'h30030070)
`define SOC_IFC_REG_CPTRA_TRNG_VALID_PAUSER                                                         (32'h70)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_PAUSER_LOCK                                                      (32'h30030074)
`define SOC_IFC_REG_CPTRA_TRNG_PAUSER_LOCK                                                          (32'h74)
`define SOC_IFC_REG_CPTRA_TRNG_PAUSER_LOCK_LOCK_LOW                                                 (0)
`define SOC_IFC_REG_CPTRA_TRNG_PAUSER_LOCK_LOCK_MASK                                                (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_0                                                           (32'h30030078)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_0                                                               (32'h78)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_1                                                           (32'h3003007c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_1                                                               (32'h7c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_2                                                           (32'h30030080)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_2                                                               (32'h80)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_3                                                           (32'h30030084)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_3                                                               (32'h84)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_4                                                           (32'h30030088)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_4                                                               (32'h88)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_5                                                           (32'h3003008c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_5                                                               (32'h8c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_6                                                           (32'h30030090)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_6                                                               (32'h90)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_7                                                           (32'h30030094)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_7                                                               (32'h94)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_8                                                           (32'h30030098)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_8                                                               (32'h98)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_9                                                           (32'h3003009c)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_9                                                               (32'h9c)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_10                                                          (32'h300300a0)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_10                                                              (32'ha0)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_DATA_11                                                          (32'h300300a4)
`define SOC_IFC_REG_CPTRA_TRNG_DATA_11                                                              (32'ha4)
`define CLP_SOC_IFC_REG_CPTRA_TRNG_STATUS                                                           (32'h300300a8)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS                                                               (32'ha8)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_REQ_LOW                                                  (0)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_REQ_MASK                                                 (32'h1)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_WR_DONE_LOW                                              (1)
`define SOC_IFC_REG_CPTRA_TRNG_STATUS_DATA_WR_DONE_MASK                                             (32'h2)
`define CLP_SOC_IFC_REG_CPTRA_FUSE_WR_DONE                                                          (32'h300300ac)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE                                                              (32'hac)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE_DONE_LOW                                                     (0)
`define SOC_IFC_REG_CPTRA_FUSE_WR_DONE_DONE_MASK                                                    (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_TIMER_CONFIG                                                          (32'h300300b0)
`define SOC_IFC_REG_CPTRA_TIMER_CONFIG                                                              (32'hb0)
`define CLP_SOC_IFC_REG_CPTRA_BOOTFSM_GO                                                            (32'h300300b4)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO                                                                (32'hb4)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO_GO_LOW                                                         (0)
`define SOC_IFC_REG_CPTRA_BOOTFSM_GO_GO_MASK                                                        (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG                                                 (32'h300300b8)
`define SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG                                                     (32'hb8)
`define CLP_SOC_IFC_REG_CPTRA_CLK_GATING_EN                                                         (32'h300300bc)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN                                                             (32'hbc)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN_CLK_GATING_EN_LOW                                           (0)
`define SOC_IFC_REG_CPTRA_CLK_GATING_EN_CLK_GATING_EN_MASK                                          (32'h1)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_0                                                 (32'h300300c0)
`define SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_0                                                     (32'hc0)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_1                                                 (32'h300300c4)
`define SOC_IFC_REG_CPTRA_GENERIC_INPUT_WIRES_1                                                     (32'hc4)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                                (32'h300300c8)
`define SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_0                                                    (32'hc8)
`define CLP_SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                                (32'h300300cc)
`define SOC_IFC_REG_CPTRA_GENERIC_OUTPUT_WIRES_1                                                    (32'hcc)
`define CLP_SOC_IFC_REG_CPTRA_HW_REV_ID                                                             (32'h300300d0)
`define SOC_IFC_REG_CPTRA_HW_REV_ID                                                                 (32'hd0)
`define CLP_SOC_IFC_REG_CPTRA_FW_REV_ID_0                                                           (32'h300300d4)
`define SOC_IFC_REG_CPTRA_FW_REV_ID_0                                                               (32'hd4)
`define CLP_SOC_IFC_REG_CPTRA_FW_REV_ID_1                                                           (32'h300300d8)
`define SOC_IFC_REG_CPTRA_FW_REV_ID_1                                                               (32'hd8)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_0                                                             (32'h30030200)
`define SOC_IFC_REG_FUSE_UDS_SEED_0                                                                 (32'h200)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_1                                                             (32'h30030204)
`define SOC_IFC_REG_FUSE_UDS_SEED_1                                                                 (32'h204)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_2                                                             (32'h30030208)
`define SOC_IFC_REG_FUSE_UDS_SEED_2                                                                 (32'h208)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_3                                                             (32'h3003020c)
`define SOC_IFC_REG_FUSE_UDS_SEED_3                                                                 (32'h20c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_4                                                             (32'h30030210)
`define SOC_IFC_REG_FUSE_UDS_SEED_4                                                                 (32'h210)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_5                                                             (32'h30030214)
`define SOC_IFC_REG_FUSE_UDS_SEED_5                                                                 (32'h214)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_6                                                             (32'h30030218)
`define SOC_IFC_REG_FUSE_UDS_SEED_6                                                                 (32'h218)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_7                                                             (32'h3003021c)
`define SOC_IFC_REG_FUSE_UDS_SEED_7                                                                 (32'h21c)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_8                                                             (32'h30030220)
`define SOC_IFC_REG_FUSE_UDS_SEED_8                                                                 (32'h220)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_9                                                             (32'h30030224)
`define SOC_IFC_REG_FUSE_UDS_SEED_9                                                                 (32'h224)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_10                                                            (32'h30030228)
`define SOC_IFC_REG_FUSE_UDS_SEED_10                                                                (32'h228)
`define CLP_SOC_IFC_REG_FUSE_UDS_SEED_11                                                            (32'h3003022c)
`define SOC_IFC_REG_FUSE_UDS_SEED_11                                                                (32'h22c)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_0                                                        (32'h30030230)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_0                                                            (32'h230)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_1                                                        (32'h30030234)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_1                                                            (32'h234)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_2                                                        (32'h30030238)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_2                                                            (32'h238)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_3                                                        (32'h3003023c)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_3                                                            (32'h23c)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_4                                                        (32'h30030240)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_4                                                            (32'h240)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_5                                                        (32'h30030244)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_5                                                            (32'h244)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_6                                                        (32'h30030248)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_6                                                            (32'h248)
`define CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_7                                                        (32'h3003024c)
`define SOC_IFC_REG_FUSE_FIELD_ENTROPY_7                                                            (32'h24c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_0                                                 (32'h30030250)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_0                                                     (32'h250)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_1                                                 (32'h30030254)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_1                                                     (32'h254)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_2                                                 (32'h30030258)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_2                                                     (32'h258)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_3                                                 (32'h3003025c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_3                                                     (32'h25c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_4                                                 (32'h30030260)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_4                                                     (32'h260)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_5                                                 (32'h30030264)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_5                                                     (32'h264)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_6                                                 (32'h30030268)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_6                                                     (32'h268)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_7                                                 (32'h3003026c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_7                                                     (32'h26c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_8                                                 (32'h30030270)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_8                                                     (32'h270)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_9                                                 (32'h30030274)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_9                                                     (32'h274)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_10                                                (32'h30030278)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_10                                                    (32'h278)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_11                                                (32'h3003027c)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_11                                                    (32'h27c)
`define CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK                                              (32'h30030280)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK                                                  (32'h280)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK_MASK_LOW                                         (0)
`define SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK_MASK_MASK                                        (32'hf)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_0                                                        (32'h30030284)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_0                                                            (32'h284)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_1                                                        (32'h30030288)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_1                                                            (32'h288)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_2                                                        (32'h3003028c)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_2                                                            (32'h28c)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_3                                                        (32'h30030290)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_3                                                            (32'h290)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_4                                                        (32'h30030294)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_4                                                            (32'h294)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_5                                                        (32'h30030298)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_5                                                            (32'h298)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_6                                                        (32'h3003029c)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_6                                                            (32'h29c)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_7                                                        (32'h300302a0)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_7                                                            (32'h2a0)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_8                                                        (32'h300302a4)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_8                                                            (32'h2a4)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_9                                                        (32'h300302a8)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_9                                                            (32'h2a8)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_10                                                       (32'h300302ac)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_10                                                           (32'h2ac)
`define CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_11                                                       (32'h300302b0)
`define SOC_IFC_REG_FUSE_OWNER_PK_HASH_11                                                           (32'h2b0)
`define CLP_SOC_IFC_REG_FUSE_FMC_KEY_MANIFEST_SVN                                                   (32'h300302b4)
`define SOC_IFC_REG_FUSE_FMC_KEY_MANIFEST_SVN                                                       (32'h2b4)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_0                                                          (32'h300302b8)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_0                                                              (32'h2b8)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_1                                                          (32'h300302bc)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_1                                                              (32'h2bc)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_2                                                          (32'h300302c0)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_2                                                              (32'h2c0)
`define CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_3                                                          (32'h300302c4)
`define SOC_IFC_REG_FUSE_RUNTIME_SVN_3                                                              (32'h2c4)
`define CLP_SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE                                                  (32'h300302c8)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE                                                      (32'h2c8)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE_DIS_LOW                                              (0)
`define SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE_DIS_MASK                                             (32'h1)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_0                                                     (32'h300302cc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_0                                                         (32'h2cc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_1                                                     (32'h300302d0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_1                                                         (32'h2d0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_2                                                     (32'h300302d4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_2                                                         (32'h2d4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_3                                                     (32'h300302d8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_3                                                         (32'h2d8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_4                                                     (32'h300302dc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_4                                                         (32'h2dc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_5                                                     (32'h300302e0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_5                                                         (32'h2e0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6                                                     (32'h300302e4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6                                                         (32'h2e4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7                                                     (32'h300302e8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7                                                         (32'h2e8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8                                                     (32'h300302ec)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8                                                         (32'h2ec)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9                                                     (32'h300302f0)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9                                                         (32'h2f0)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10                                                    (32'h300302f4)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10                                                        (32'h2f4)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_11                                                    (32'h300302f8)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_11                                                        (32'h2f8)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_12                                                    (32'h300302fc)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_12                                                        (32'h2fc)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_13                                                    (32'h30030300)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_13                                                        (32'h300)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_14                                                    (32'h30030304)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_14                                                        (32'h304)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_15                                                    (32'h30030308)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_15                                                        (32'h308)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_16                                                    (32'h3003030c)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_16                                                        (32'h30c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_17                                                    (32'h30030310)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_17                                                        (32'h310)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_18                                                    (32'h30030314)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_18                                                        (32'h314)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_19                                                    (32'h30030318)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_19                                                        (32'h318)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_20                                                    (32'h3003031c)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_20                                                        (32'h31c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_21                                                    (32'h30030320)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_21                                                        (32'h320)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_22                                                    (32'h30030324)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_22                                                        (32'h324)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_23                                                    (32'h30030328)
`define SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_23                                                        (32'h328)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                                  (32'h3003032c)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_0                                                      (32'h32c)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                                  (32'h30030330)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_1                                                      (32'h330)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                                  (32'h30030334)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_2                                                      (32'h334)
`define CLP_SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                                  (32'h30030338)
`define SOC_IFC_REG_FUSE_IDEVID_MANUF_HSM_ID_3                                                      (32'h338)
`define CLP_SOC_IFC_REG_FUSE_LIFE_CYCLE                                                             (32'h3003033c)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE                                                                 (32'h33c)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE_LIFE_CYCLE_LOW                                                  (0)
`define SOC_IFC_REG_FUSE_LIFE_CYCLE_LIFE_CYCLE_MASK                                                 (32'h3)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_0                                                          (32'h30030600)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_0                                                              (32'h600)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_1                                                          (32'h30030604)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_1                                                              (32'h604)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_2                                                          (32'h30030608)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_2                                                              (32'h608)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_3                                                          (32'h3003060c)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_3                                                              (32'h60c)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_4                                                          (32'h30030610)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_4                                                              (32'h610)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_5                                                          (32'h30030614)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_5                                                              (32'h614)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_6                                                          (32'h30030618)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_6                                                              (32'h618)
`define CLP_SOC_IFC_REG_INTERNAL_OBF_KEY_7                                                          (32'h3003061c)
`define SOC_IFC_REG_INTERNAL_OBF_KEY_7                                                              (32'h61c)
`define CLP_SOC_IFC_REG_INTERNAL_ICCM_LOCK                                                          (32'h30030620)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK                                                              (32'h620)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK_LOCK_LOW                                                     (0)
`define SOC_IFC_REG_INTERNAL_ICCM_LOCK_LOCK_MASK                                                    (32'h1)
`define CLP_SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET                                                    (32'h30030624)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET                                                        (32'h624)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_CORE_RST_LOW                                           (0)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_CORE_RST_MASK                                          (32'h1)
`define CLP_SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES                                        (32'h30030628)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES                                            (32'h628)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES_WAIT_CYCLES_LOW                            (0)
`define SOC_IFC_REG_INTERNAL_FW_UPDATE_RESET_WAIT_CYCLES_WAIT_CYCLES_MASK                           (32'hff)
`define CLP_SOC_IFC_REG_INTERNAL_NMI_VECTOR                                                         (32'h3003062c)
`define SOC_IFC_REG_INTERNAL_NMI_VECTOR                                                             (32'h62c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_START                                                         (32'h30030800)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                              (32'h30030800)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R                                                  (32'h800)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_LOW                                     (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_ERROR_EN_MASK                                    (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_LOW                                     (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_GLOBAL_INTR_EN_R_NOTIF_EN_MASK                                    (32'h2)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                               (32'h30030804)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R                                                   (32'h804)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_LOW                             (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INTERNAL_EN_MASK                            (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INV_DEV_EN_LOW                              (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_INV_DEV_EN_MASK                             (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_CMD_FAIL_EN_LOW                             (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_CMD_FAIL_EN_MASK                            (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_BAD_FUSE_EN_LOW                             (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_BAD_FUSE_EN_MASK                            (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_ICCM_BLOCKED_EN_LOW                         (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_ICCM_BLOCKED_EN_MASK                        (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_MBOX_ECC_UNC_EN_LOW                         (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_EN_R_ERROR_MBOX_ECC_UNC_EN_MASK                        (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                               (32'h30030808)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R                                                   (32'h808)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_AVAIL_EN_LOW                            (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_CMD_AVAIL_EN_MASK                           (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_MBOX_ECC_COR_EN_LOW                         (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_MBOX_ECC_COR_EN_MASK                        (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_DEBUG_LOCKED_EN_LOW                         (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_EN_R_NOTIF_DEBUG_LOCKED_EN_MASK                        (32'h4)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                           (32'h3003080c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R                                               (32'h80c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_LOW                                   (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_GLOBAL_INTR_R_AGG_STS_MASK                                  (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                           (32'h30030810)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R                                               (32'h810)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_LOW                                   (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_GLOBAL_INTR_R_AGG_STS_MASK                                  (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                         (32'h30030814)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R                                             (32'h814)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_LOW                      (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INTERNAL_STS_MASK                     (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INV_DEV_STS_LOW                       (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_INV_DEV_STS_MASK                      (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_CMD_FAIL_STS_LOW                      (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_CMD_FAIL_STS_MASK                     (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_BAD_FUSE_STS_LOW                      (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_BAD_FUSE_STS_MASK                     (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_ICCM_BLOCKED_STS_LOW                  (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_ICCM_BLOCKED_STS_MASK                 (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_MBOX_ECC_UNC_STS_LOW                  (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_R_ERROR_MBOX_ECC_UNC_STS_MASK                 (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                         (32'h30030818)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R                                             (32'h818)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_AVAIL_STS_LOW                     (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_CMD_AVAIL_STS_MASK                    (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_MBOX_ECC_COR_STS_LOW                  (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_MBOX_ECC_COR_STS_MASK                 (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_DEBUG_LOCKED_STS_LOW                  (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTERNAL_INTR_R_NOTIF_DEBUG_LOCKED_STS_MASK                 (32'h4)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                             (32'h3003081c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R                                                 (32'h81c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_LOW                         (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INTERNAL_TRIG_MASK                        (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INV_DEV_TRIG_LOW                          (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_INV_DEV_TRIG_MASK                         (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_CMD_FAIL_TRIG_LOW                         (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_CMD_FAIL_TRIG_MASK                        (32'h4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_BAD_FUSE_TRIG_LOW                         (3)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_BAD_FUSE_TRIG_MASK                        (32'h8)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_ICCM_BLOCKED_TRIG_LOW                     (4)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_ICCM_BLOCKED_TRIG_MASK                    (32'h10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_MBOX_ECC_UNC_TRIG_LOW                     (5)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTR_TRIG_R_ERROR_MBOX_ECC_UNC_TRIG_MASK                    (32'h20)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                             (32'h30030820)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R                                                 (32'h820)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_AVAIL_TRIG_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_CMD_AVAIL_TRIG_MASK                       (32'h1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_MBOX_ECC_COR_TRIG_LOW                     (1)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_MBOX_ECC_COR_TRIG_MASK                    (32'h2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_DEBUG_LOCKED_TRIG_LOW                     (2)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_INTR_TRIG_R_NOTIF_DEBUG_LOCKED_TRIG_MASK                    (32'h4)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                   (32'h30030900)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_R                                       (32'h900)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_R                                    (32'h30030904)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_R                                        (32'h904)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_R                                   (32'h30030908)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_R                                       (32'h908)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_R                                   (32'h3003090c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_R                                       (32'h90c)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_R                               (32'h30030910)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_R                                   (32'h910)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_R                               (32'h30030914)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_R                                   (32'h914)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_R                                  (32'h30030980)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_R                                      (32'h980)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_R                               (32'h30030984)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_R                                   (32'h984)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                               (32'h30030988)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_R                                   (32'h988)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                              (32'h30030a00)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R                                  (32'ha00)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INTERNAL_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R                               (32'h30030a04)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R                                   (32'ha04)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R_PULSE_LOW                         (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_INV_DEV_INTR_COUNT_INCR_R_PULSE_MASK                        (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R                              (32'h30030a08)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R                                  (32'ha08)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_CMD_FAIL_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R                              (32'h30030a0c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R                                  (32'ha0c)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R_PULSE_LOW                        (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_BAD_FUSE_INTR_COUNT_INCR_R_PULSE_MASK                       (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R                          (32'h30030a10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R                              (32'ha10)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_ICCM_BLOCKED_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R                          (32'h30030a14)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R                              (32'ha14)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_ERROR_MBOX_ECC_UNC_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R                             (32'h30030a18)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R                                 (32'ha18)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R_PULSE_LOW                       (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_CMD_AVAIL_INTR_COUNT_INCR_R_PULSE_MASK                      (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R                          (32'h30030a1c)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R                              (32'ha1c)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_MBOX_ECC_COR_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)
`define CLP_SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                          (32'h30030a20)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R                              (32'ha20)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R_PULSE_LOW                    (0)
`define SOC_IFC_REG_INTR_BLOCK_RF_NOTIF_DEBUG_LOCKED_INTR_COUNT_INCR_R_PULSE_MASK                   (32'h1)


`endif